magic
tech sky130A
magscale 1 2
timestamp 1617639612
<< obsli1 >>
rect 43545 2533 512963 700995
<< obsm1 >>
rect 566 1980 582820 701808
<< metal2 >>
rect 7074 703520 7186 704960
rect 21242 703520 21354 704960
rect 35502 703520 35614 704960
rect 49762 703520 49874 704960
rect 64022 703520 64134 704960
rect 78282 703520 78394 704960
rect 92450 703520 92562 704960
rect 106710 703520 106822 704960
rect 120970 703520 121082 704960
rect 135230 703520 135342 704960
rect 149490 703520 149602 704960
rect 163750 703520 163862 704960
rect 177918 703520 178030 704960
rect 192178 703520 192290 704960
rect 206438 703520 206550 704960
rect 220698 703520 220810 704960
rect 234958 703520 235070 704960
rect 249218 703520 249330 704960
rect 263386 703520 263498 704960
rect 277646 703520 277758 704960
rect 291906 703520 292018 704960
rect 306166 703520 306278 704960
rect 320426 703520 320538 704960
rect 334686 703520 334798 704960
rect 348854 703520 348966 704960
rect 363114 703520 363226 704960
rect 377374 703520 377486 704960
rect 391634 703520 391746 704960
rect 405894 703520 406006 704960
rect 420154 703520 420266 704960
rect 434322 703520 434434 704960
rect 448582 703520 448694 704960
rect 462842 703520 462954 704960
rect 477102 703520 477214 704960
rect 491362 703520 491474 704960
rect 505622 703520 505734 704960
rect 519790 703520 519902 704960
rect 534050 703520 534162 704960
rect 548310 703520 548422 704960
rect 562570 703520 562682 704960
rect 576830 703520 576942 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6338 -960 6450 480
rect 7534 -960 7646 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11030 -960 11142 480
rect 12226 -960 12338 480
rect 13422 -960 13534 480
rect 14618 -960 14730 480
rect 15814 -960 15926 480
rect 16918 -960 17030 480
rect 18114 -960 18226 480
rect 19310 -960 19422 480
rect 20506 -960 20618 480
rect 21610 -960 21722 480
rect 22806 -960 22918 480
rect 24002 -960 24114 480
rect 25198 -960 25310 480
rect 26302 -960 26414 480
rect 27498 -960 27610 480
rect 28694 -960 28806 480
rect 29890 -960 30002 480
rect 31086 -960 31198 480
rect 32190 -960 32302 480
rect 33386 -960 33498 480
rect 34582 -960 34694 480
rect 35778 -960 35890 480
rect 36882 -960 36994 480
rect 38078 -960 38190 480
rect 39274 -960 39386 480
rect 40470 -960 40582 480
rect 41666 -960 41778 480
rect 42770 -960 42882 480
rect 43966 -960 44078 480
rect 45162 -960 45274 480
rect 46358 -960 46470 480
rect 47462 -960 47574 480
rect 48658 -960 48770 480
rect 49854 -960 49966 480
rect 51050 -960 51162 480
rect 52154 -960 52266 480
rect 53350 -960 53462 480
rect 54546 -960 54658 480
rect 55742 -960 55854 480
rect 56938 -960 57050 480
rect 58042 -960 58154 480
rect 59238 -960 59350 480
rect 60434 -960 60546 480
rect 61630 -960 61742 480
rect 62734 -960 62846 480
rect 63930 -960 64042 480
rect 65126 -960 65238 480
rect 66322 -960 66434 480
rect 67518 -960 67630 480
rect 68622 -960 68734 480
rect 69818 -960 69930 480
rect 71014 -960 71126 480
rect 72210 -960 72322 480
rect 73314 -960 73426 480
rect 74510 -960 74622 480
rect 75706 -960 75818 480
rect 76902 -960 77014 480
rect 78006 -960 78118 480
rect 79202 -960 79314 480
rect 80398 -960 80510 480
rect 81594 -960 81706 480
rect 82790 -960 82902 480
rect 83894 -960 84006 480
rect 85090 -960 85202 480
rect 86286 -960 86398 480
rect 87482 -960 87594 480
rect 88586 -960 88698 480
rect 89782 -960 89894 480
rect 90978 -960 91090 480
rect 92174 -960 92286 480
rect 93370 -960 93482 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99166 -960 99278 480
rect 100362 -960 100474 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103858 -960 103970 480
rect 105054 -960 105166 480
rect 106250 -960 106362 480
rect 107446 -960 107558 480
rect 108642 -960 108754 480
rect 109746 -960 109858 480
rect 110942 -960 111054 480
rect 112138 -960 112250 480
rect 113334 -960 113446 480
rect 114438 -960 114550 480
rect 115634 -960 115746 480
rect 116830 -960 116942 480
rect 118026 -960 118138 480
rect 119222 -960 119334 480
rect 120326 -960 120438 480
rect 121522 -960 121634 480
rect 122718 -960 122830 480
rect 123914 -960 124026 480
rect 125018 -960 125130 480
rect 126214 -960 126326 480
rect 127410 -960 127522 480
rect 128606 -960 128718 480
rect 129710 -960 129822 480
rect 130906 -960 131018 480
rect 132102 -960 132214 480
rect 133298 -960 133410 480
rect 134494 -960 134606 480
rect 135598 -960 135710 480
rect 136794 -960 136906 480
rect 137990 -960 138102 480
rect 139186 -960 139298 480
rect 140290 -960 140402 480
rect 141486 -960 141598 480
rect 142682 -960 142794 480
rect 143878 -960 143990 480
rect 145074 -960 145186 480
rect 146178 -960 146290 480
rect 147374 -960 147486 480
rect 148570 -960 148682 480
rect 149766 -960 149878 480
rect 150870 -960 150982 480
rect 152066 -960 152178 480
rect 153262 -960 153374 480
rect 154458 -960 154570 480
rect 155562 -960 155674 480
rect 156758 -960 156870 480
rect 157954 -960 158066 480
rect 159150 -960 159262 480
rect 160346 -960 160458 480
rect 161450 -960 161562 480
rect 162646 -960 162758 480
rect 163842 -960 163954 480
rect 165038 -960 165150 480
rect 166142 -960 166254 480
rect 167338 -960 167450 480
rect 168534 -960 168646 480
rect 169730 -960 169842 480
rect 170926 -960 171038 480
rect 172030 -960 172142 480
rect 173226 -960 173338 480
rect 174422 -960 174534 480
rect 175618 -960 175730 480
rect 176722 -960 176834 480
rect 177918 -960 178030 480
rect 179114 -960 179226 480
rect 180310 -960 180422 480
rect 181414 -960 181526 480
rect 182610 -960 182722 480
rect 183806 -960 183918 480
rect 185002 -960 185114 480
rect 186198 -960 186310 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190890 -960 191002 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202574 -960 202686 480
rect 203770 -960 203882 480
rect 204966 -960 205078 480
rect 206162 -960 206274 480
rect 207266 -960 207378 480
rect 208462 -960 208574 480
rect 209658 -960 209770 480
rect 210854 -960 210966 480
rect 212050 -960 212162 480
rect 213154 -960 213266 480
rect 214350 -960 214462 480
rect 215546 -960 215658 480
rect 216742 -960 216854 480
rect 217846 -960 217958 480
rect 219042 -960 219154 480
rect 220238 -960 220350 480
rect 221434 -960 221546 480
rect 222630 -960 222742 480
rect 223734 -960 223846 480
rect 224930 -960 225042 480
rect 226126 -960 226238 480
rect 227322 -960 227434 480
rect 228426 -960 228538 480
rect 229622 -960 229734 480
rect 230818 -960 230930 480
rect 232014 -960 232126 480
rect 233118 -960 233230 480
rect 234314 -960 234426 480
rect 235510 -960 235622 480
rect 236706 -960 236818 480
rect 237902 -960 238014 480
rect 239006 -960 239118 480
rect 240202 -960 240314 480
rect 241398 -960 241510 480
rect 242594 -960 242706 480
rect 243698 -960 243810 480
rect 244894 -960 245006 480
rect 246090 -960 246202 480
rect 247286 -960 247398 480
rect 248482 -960 248594 480
rect 249586 -960 249698 480
rect 250782 -960 250894 480
rect 251978 -960 252090 480
rect 253174 -960 253286 480
rect 254278 -960 254390 480
rect 255474 -960 255586 480
rect 256670 -960 256782 480
rect 257866 -960 257978 480
rect 258970 -960 259082 480
rect 260166 -960 260278 480
rect 261362 -960 261474 480
rect 262558 -960 262670 480
rect 263754 -960 263866 480
rect 264858 -960 264970 480
rect 266054 -960 266166 480
rect 267250 -960 267362 480
rect 268446 -960 268558 480
rect 269550 -960 269662 480
rect 270746 -960 270858 480
rect 271942 -960 272054 480
rect 273138 -960 273250 480
rect 274334 -960 274446 480
rect 275438 -960 275550 480
rect 276634 -960 276746 480
rect 277830 -960 277942 480
rect 279026 -960 279138 480
rect 280130 -960 280242 480
rect 281326 -960 281438 480
rect 282522 -960 282634 480
rect 283718 -960 283830 480
rect 284822 -960 284934 480
rect 286018 -960 286130 480
rect 287214 -960 287326 480
rect 288410 -960 288522 480
rect 289606 -960 289718 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295402 -960 295514 480
rect 296598 -960 296710 480
rect 297794 -960 297906 480
rect 298990 -960 299102 480
rect 300186 -960 300298 480
rect 301290 -960 301402 480
rect 302486 -960 302598 480
rect 303682 -960 303794 480
rect 304878 -960 304990 480
rect 305982 -960 306094 480
rect 307178 -960 307290 480
rect 308374 -960 308486 480
rect 309570 -960 309682 480
rect 310674 -960 310786 480
rect 311870 -960 311982 480
rect 313066 -960 313178 480
rect 314262 -960 314374 480
rect 315458 -960 315570 480
rect 316562 -960 316674 480
rect 317758 -960 317870 480
rect 318954 -960 319066 480
rect 320150 -960 320262 480
rect 321254 -960 321366 480
rect 322450 -960 322562 480
rect 323646 -960 323758 480
rect 324842 -960 324954 480
rect 326038 -960 326150 480
rect 327142 -960 327254 480
rect 328338 -960 328450 480
rect 329534 -960 329646 480
rect 330730 -960 330842 480
rect 331834 -960 331946 480
rect 333030 -960 333142 480
rect 334226 -960 334338 480
rect 335422 -960 335534 480
rect 336526 -960 336638 480
rect 337722 -960 337834 480
rect 338918 -960 339030 480
rect 340114 -960 340226 480
rect 341310 -960 341422 480
rect 342414 -960 342526 480
rect 343610 -960 343722 480
rect 344806 -960 344918 480
rect 346002 -960 346114 480
rect 347106 -960 347218 480
rect 348302 -960 348414 480
rect 349498 -960 349610 480
rect 350694 -960 350806 480
rect 351890 -960 352002 480
rect 352994 -960 353106 480
rect 354190 -960 354302 480
rect 355386 -960 355498 480
rect 356582 -960 356694 480
rect 357686 -960 357798 480
rect 358882 -960 358994 480
rect 360078 -960 360190 480
rect 361274 -960 361386 480
rect 362378 -960 362490 480
rect 363574 -960 363686 480
rect 364770 -960 364882 480
rect 365966 -960 366078 480
rect 367162 -960 367274 480
rect 368266 -960 368378 480
rect 369462 -960 369574 480
rect 370658 -960 370770 480
rect 371854 -960 371966 480
rect 372958 -960 373070 480
rect 374154 -960 374266 480
rect 375350 -960 375462 480
rect 376546 -960 376658 480
rect 377742 -960 377854 480
rect 378846 -960 378958 480
rect 380042 -960 380154 480
rect 381238 -960 381350 480
rect 382434 -960 382546 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394118 -960 394230 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398810 -960 398922 480
rect 400006 -960 400118 480
rect 401202 -960 401314 480
rect 402398 -960 402510 480
rect 403594 -960 403706 480
rect 404698 -960 404810 480
rect 405894 -960 406006 480
rect 407090 -960 407202 480
rect 408286 -960 408398 480
rect 409390 -960 409502 480
rect 410586 -960 410698 480
rect 411782 -960 411894 480
rect 412978 -960 413090 480
rect 414082 -960 414194 480
rect 415278 -960 415390 480
rect 416474 -960 416586 480
rect 417670 -960 417782 480
rect 418866 -960 418978 480
rect 419970 -960 420082 480
rect 421166 -960 421278 480
rect 422362 -960 422474 480
rect 423558 -960 423670 480
rect 424662 -960 424774 480
rect 425858 -960 425970 480
rect 427054 -960 427166 480
rect 428250 -960 428362 480
rect 429446 -960 429558 480
rect 430550 -960 430662 480
rect 431746 -960 431858 480
rect 432942 -960 433054 480
rect 434138 -960 434250 480
rect 435242 -960 435354 480
rect 436438 -960 436550 480
rect 437634 -960 437746 480
rect 438830 -960 438942 480
rect 439934 -960 440046 480
rect 441130 -960 441242 480
rect 442326 -960 442438 480
rect 443522 -960 443634 480
rect 444718 -960 444830 480
rect 445822 -960 445934 480
rect 447018 -960 447130 480
rect 448214 -960 448326 480
rect 449410 -960 449522 480
rect 450514 -960 450626 480
rect 451710 -960 451822 480
rect 452906 -960 453018 480
rect 454102 -960 454214 480
rect 455298 -960 455410 480
rect 456402 -960 456514 480
rect 457598 -960 457710 480
rect 458794 -960 458906 480
rect 459990 -960 460102 480
rect 461094 -960 461206 480
rect 462290 -960 462402 480
rect 463486 -960 463598 480
rect 464682 -960 464794 480
rect 465786 -960 465898 480
rect 466982 -960 467094 480
rect 468178 -960 468290 480
rect 469374 -960 469486 480
rect 470570 -960 470682 480
rect 471674 -960 471786 480
rect 472870 -960 472982 480
rect 474066 -960 474178 480
rect 475262 -960 475374 480
rect 476366 -960 476478 480
rect 477562 -960 477674 480
rect 478758 -960 478870 480
rect 479954 -960 480066 480
rect 481150 -960 481262 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484646 -960 484758 480
rect 485842 -960 485954 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491638 -960 491750 480
rect 492834 -960 492946 480
rect 494030 -960 494142 480
rect 495226 -960 495338 480
rect 496422 -960 496534 480
rect 497526 -960 497638 480
rect 498722 -960 498834 480
rect 499918 -960 500030 480
rect 501114 -960 501226 480
rect 502218 -960 502330 480
rect 503414 -960 503526 480
rect 504610 -960 504722 480
rect 505806 -960 505918 480
rect 507002 -960 507114 480
rect 508106 -960 508218 480
rect 509302 -960 509414 480
rect 510498 -960 510610 480
rect 511694 -960 511806 480
rect 512798 -960 512910 480
rect 513994 -960 514106 480
rect 515190 -960 515302 480
rect 516386 -960 516498 480
rect 517490 -960 517602 480
rect 518686 -960 518798 480
rect 519882 -960 519994 480
rect 521078 -960 521190 480
rect 522274 -960 522386 480
rect 523378 -960 523490 480
rect 524574 -960 524686 480
rect 525770 -960 525882 480
rect 526966 -960 527078 480
rect 528070 -960 528182 480
rect 529266 -960 529378 480
rect 530462 -960 530574 480
rect 531658 -960 531770 480
rect 532854 -960 532966 480
rect 533958 -960 534070 480
rect 535154 -960 535266 480
rect 536350 -960 536462 480
rect 537546 -960 537658 480
rect 538650 -960 538762 480
rect 539846 -960 539958 480
rect 541042 -960 541154 480
rect 542238 -960 542350 480
rect 543342 -960 543454 480
rect 544538 -960 544650 480
rect 545734 -960 545846 480
rect 546930 -960 547042 480
rect 548126 -960 548238 480
rect 549230 -960 549342 480
rect 550426 -960 550538 480
rect 551622 -960 551734 480
rect 552818 -960 552930 480
rect 553922 -960 554034 480
rect 555118 -960 555230 480
rect 556314 -960 556426 480
rect 557510 -960 557622 480
rect 558706 -960 558818 480
rect 559810 -960 559922 480
rect 561006 -960 561118 480
rect 562202 -960 562314 480
rect 563398 -960 563510 480
rect 564502 -960 564614 480
rect 565698 -960 565810 480
rect 566894 -960 567006 480
rect 568090 -960 568202 480
rect 569194 -960 569306 480
rect 570390 -960 570502 480
rect 571586 -960 571698 480
rect 572782 -960 572894 480
rect 573978 -960 574090 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577474 -960 577586 480
rect 578670 -960 578782 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 7018 703520
rect 7242 703464 21186 703520
rect 21410 703464 35446 703520
rect 35670 703464 49706 703520
rect 49930 703464 63966 703520
rect 64190 703464 78226 703520
rect 78450 703464 92394 703520
rect 92618 703464 106654 703520
rect 106878 703464 120914 703520
rect 121138 703464 135174 703520
rect 135398 703464 149434 703520
rect 149658 703464 163694 703520
rect 163918 703464 177862 703520
rect 178086 703464 192122 703520
rect 192346 703464 206382 703520
rect 206606 703464 220642 703520
rect 220866 703464 234902 703520
rect 235126 703464 249162 703520
rect 249386 703464 263330 703520
rect 263554 703464 277590 703520
rect 277814 703464 291850 703520
rect 292074 703464 306110 703520
rect 306334 703464 320370 703520
rect 320594 703464 334630 703520
rect 334854 703464 348798 703520
rect 349022 703464 363058 703520
rect 363282 703464 377318 703520
rect 377542 703464 391578 703520
rect 391802 703464 405838 703520
rect 406062 703464 420098 703520
rect 420322 703464 434266 703520
rect 434490 703464 448526 703520
rect 448750 703464 462786 703520
rect 463010 703464 477046 703520
rect 477270 703464 491306 703520
rect 491530 703464 505566 703520
rect 505790 703464 519734 703520
rect 519958 703464 533994 703520
rect 534218 703464 548254 703520
rect 548478 703464 562514 703520
rect 562738 703464 576774 703520
rect 576998 703464 583432 703520
rect 572 536 583432 703464
rect 710 480 1590 536
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6282 536
rect 6506 480 7478 536
rect 7702 480 8674 536
rect 8898 480 9870 536
rect 10094 480 10974 536
rect 11198 480 12170 536
rect 12394 480 13366 536
rect 13590 480 14562 536
rect 14786 480 15758 536
rect 15982 480 16862 536
rect 17086 480 18058 536
rect 18282 480 19254 536
rect 19478 480 20450 536
rect 20674 480 21554 536
rect 21778 480 22750 536
rect 22974 480 23946 536
rect 24170 480 25142 536
rect 25366 480 26246 536
rect 26470 480 27442 536
rect 27666 480 28638 536
rect 28862 480 29834 536
rect 30058 480 31030 536
rect 31254 480 32134 536
rect 32358 480 33330 536
rect 33554 480 34526 536
rect 34750 480 35722 536
rect 35946 480 36826 536
rect 37050 480 38022 536
rect 38246 480 39218 536
rect 39442 480 40414 536
rect 40638 480 41610 536
rect 41834 480 42714 536
rect 42938 480 43910 536
rect 44134 480 45106 536
rect 45330 480 46302 536
rect 46526 480 47406 536
rect 47630 480 48602 536
rect 48826 480 49798 536
rect 50022 480 50994 536
rect 51218 480 52098 536
rect 52322 480 53294 536
rect 53518 480 54490 536
rect 54714 480 55686 536
rect 55910 480 56882 536
rect 57106 480 57986 536
rect 58210 480 59182 536
rect 59406 480 60378 536
rect 60602 480 61574 536
rect 61798 480 62678 536
rect 62902 480 63874 536
rect 64098 480 65070 536
rect 65294 480 66266 536
rect 66490 480 67462 536
rect 67686 480 68566 536
rect 68790 480 69762 536
rect 69986 480 70958 536
rect 71182 480 72154 536
rect 72378 480 73258 536
rect 73482 480 74454 536
rect 74678 480 75650 536
rect 75874 480 76846 536
rect 77070 480 77950 536
rect 78174 480 79146 536
rect 79370 480 80342 536
rect 80566 480 81538 536
rect 81762 480 82734 536
rect 82958 480 83838 536
rect 84062 480 85034 536
rect 85258 480 86230 536
rect 86454 480 87426 536
rect 87650 480 88530 536
rect 88754 480 89726 536
rect 89950 480 90922 536
rect 91146 480 92118 536
rect 92342 480 93314 536
rect 93538 480 94418 536
rect 94642 480 95614 536
rect 95838 480 96810 536
rect 97034 480 98006 536
rect 98230 480 99110 536
rect 99334 480 100306 536
rect 100530 480 101502 536
rect 101726 480 102698 536
rect 102922 480 103802 536
rect 104026 480 104998 536
rect 105222 480 106194 536
rect 106418 480 107390 536
rect 107614 480 108586 536
rect 108810 480 109690 536
rect 109914 480 110886 536
rect 111110 480 112082 536
rect 112306 480 113278 536
rect 113502 480 114382 536
rect 114606 480 115578 536
rect 115802 480 116774 536
rect 116998 480 117970 536
rect 118194 480 119166 536
rect 119390 480 120270 536
rect 120494 480 121466 536
rect 121690 480 122662 536
rect 122886 480 123858 536
rect 124082 480 124962 536
rect 125186 480 126158 536
rect 126382 480 127354 536
rect 127578 480 128550 536
rect 128774 480 129654 536
rect 129878 480 130850 536
rect 131074 480 132046 536
rect 132270 480 133242 536
rect 133466 480 134438 536
rect 134662 480 135542 536
rect 135766 480 136738 536
rect 136962 480 137934 536
rect 138158 480 139130 536
rect 139354 480 140234 536
rect 140458 480 141430 536
rect 141654 480 142626 536
rect 142850 480 143822 536
rect 144046 480 145018 536
rect 145242 480 146122 536
rect 146346 480 147318 536
rect 147542 480 148514 536
rect 148738 480 149710 536
rect 149934 480 150814 536
rect 151038 480 152010 536
rect 152234 480 153206 536
rect 153430 480 154402 536
rect 154626 480 155506 536
rect 155730 480 156702 536
rect 156926 480 157898 536
rect 158122 480 159094 536
rect 159318 480 160290 536
rect 160514 480 161394 536
rect 161618 480 162590 536
rect 162814 480 163786 536
rect 164010 480 164982 536
rect 165206 480 166086 536
rect 166310 480 167282 536
rect 167506 480 168478 536
rect 168702 480 169674 536
rect 169898 480 170870 536
rect 171094 480 171974 536
rect 172198 480 173170 536
rect 173394 480 174366 536
rect 174590 480 175562 536
rect 175786 480 176666 536
rect 176890 480 177862 536
rect 178086 480 179058 536
rect 179282 480 180254 536
rect 180478 480 181358 536
rect 181582 480 182554 536
rect 182778 480 183750 536
rect 183974 480 184946 536
rect 185170 480 186142 536
rect 186366 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190834 536
rect 191058 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202518 536
rect 202742 480 203714 536
rect 203938 480 204910 536
rect 205134 480 206106 536
rect 206330 480 207210 536
rect 207434 480 208406 536
rect 208630 480 209602 536
rect 209826 480 210798 536
rect 211022 480 211994 536
rect 212218 480 213098 536
rect 213322 480 214294 536
rect 214518 480 215490 536
rect 215714 480 216686 536
rect 216910 480 217790 536
rect 218014 480 218986 536
rect 219210 480 220182 536
rect 220406 480 221378 536
rect 221602 480 222574 536
rect 222798 480 223678 536
rect 223902 480 224874 536
rect 225098 480 226070 536
rect 226294 480 227266 536
rect 227490 480 228370 536
rect 228594 480 229566 536
rect 229790 480 230762 536
rect 230986 480 231958 536
rect 232182 480 233062 536
rect 233286 480 234258 536
rect 234482 480 235454 536
rect 235678 480 236650 536
rect 236874 480 237846 536
rect 238070 480 238950 536
rect 239174 480 240146 536
rect 240370 480 241342 536
rect 241566 480 242538 536
rect 242762 480 243642 536
rect 243866 480 244838 536
rect 245062 480 246034 536
rect 246258 480 247230 536
rect 247454 480 248426 536
rect 248650 480 249530 536
rect 249754 480 250726 536
rect 250950 480 251922 536
rect 252146 480 253118 536
rect 253342 480 254222 536
rect 254446 480 255418 536
rect 255642 480 256614 536
rect 256838 480 257810 536
rect 258034 480 258914 536
rect 259138 480 260110 536
rect 260334 480 261306 536
rect 261530 480 262502 536
rect 262726 480 263698 536
rect 263922 480 264802 536
rect 265026 480 265998 536
rect 266222 480 267194 536
rect 267418 480 268390 536
rect 268614 480 269494 536
rect 269718 480 270690 536
rect 270914 480 271886 536
rect 272110 480 273082 536
rect 273306 480 274278 536
rect 274502 480 275382 536
rect 275606 480 276578 536
rect 276802 480 277774 536
rect 277998 480 278970 536
rect 279194 480 280074 536
rect 280298 480 281270 536
rect 281494 480 282466 536
rect 282690 480 283662 536
rect 283886 480 284766 536
rect 284990 480 285962 536
rect 286186 480 287158 536
rect 287382 480 288354 536
rect 288578 480 289550 536
rect 289774 480 290654 536
rect 290878 480 291850 536
rect 292074 480 293046 536
rect 293270 480 294242 536
rect 294466 480 295346 536
rect 295570 480 296542 536
rect 296766 480 297738 536
rect 297962 480 298934 536
rect 299158 480 300130 536
rect 300354 480 301234 536
rect 301458 480 302430 536
rect 302654 480 303626 536
rect 303850 480 304822 536
rect 305046 480 305926 536
rect 306150 480 307122 536
rect 307346 480 308318 536
rect 308542 480 309514 536
rect 309738 480 310618 536
rect 310842 480 311814 536
rect 312038 480 313010 536
rect 313234 480 314206 536
rect 314430 480 315402 536
rect 315626 480 316506 536
rect 316730 480 317702 536
rect 317926 480 318898 536
rect 319122 480 320094 536
rect 320318 480 321198 536
rect 321422 480 322394 536
rect 322618 480 323590 536
rect 323814 480 324786 536
rect 325010 480 325982 536
rect 326206 480 327086 536
rect 327310 480 328282 536
rect 328506 480 329478 536
rect 329702 480 330674 536
rect 330898 480 331778 536
rect 332002 480 332974 536
rect 333198 480 334170 536
rect 334394 480 335366 536
rect 335590 480 336470 536
rect 336694 480 337666 536
rect 337890 480 338862 536
rect 339086 480 340058 536
rect 340282 480 341254 536
rect 341478 480 342358 536
rect 342582 480 343554 536
rect 343778 480 344750 536
rect 344974 480 345946 536
rect 346170 480 347050 536
rect 347274 480 348246 536
rect 348470 480 349442 536
rect 349666 480 350638 536
rect 350862 480 351834 536
rect 352058 480 352938 536
rect 353162 480 354134 536
rect 354358 480 355330 536
rect 355554 480 356526 536
rect 356750 480 357630 536
rect 357854 480 358826 536
rect 359050 480 360022 536
rect 360246 480 361218 536
rect 361442 480 362322 536
rect 362546 480 363518 536
rect 363742 480 364714 536
rect 364938 480 365910 536
rect 366134 480 367106 536
rect 367330 480 368210 536
rect 368434 480 369406 536
rect 369630 480 370602 536
rect 370826 480 371798 536
rect 372022 480 372902 536
rect 373126 480 374098 536
rect 374322 480 375294 536
rect 375518 480 376490 536
rect 376714 480 377686 536
rect 377910 480 378790 536
rect 379014 480 379986 536
rect 380210 480 381182 536
rect 381406 480 382378 536
rect 382602 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394062 536
rect 394286 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398754 536
rect 398978 480 399950 536
rect 400174 480 401146 536
rect 401370 480 402342 536
rect 402566 480 403538 536
rect 403762 480 404642 536
rect 404866 480 405838 536
rect 406062 480 407034 536
rect 407258 480 408230 536
rect 408454 480 409334 536
rect 409558 480 410530 536
rect 410754 480 411726 536
rect 411950 480 412922 536
rect 413146 480 414026 536
rect 414250 480 415222 536
rect 415446 480 416418 536
rect 416642 480 417614 536
rect 417838 480 418810 536
rect 419034 480 419914 536
rect 420138 480 421110 536
rect 421334 480 422306 536
rect 422530 480 423502 536
rect 423726 480 424606 536
rect 424830 480 425802 536
rect 426026 480 426998 536
rect 427222 480 428194 536
rect 428418 480 429390 536
rect 429614 480 430494 536
rect 430718 480 431690 536
rect 431914 480 432886 536
rect 433110 480 434082 536
rect 434306 480 435186 536
rect 435410 480 436382 536
rect 436606 480 437578 536
rect 437802 480 438774 536
rect 438998 480 439878 536
rect 440102 480 441074 536
rect 441298 480 442270 536
rect 442494 480 443466 536
rect 443690 480 444662 536
rect 444886 480 445766 536
rect 445990 480 446962 536
rect 447186 480 448158 536
rect 448382 480 449354 536
rect 449578 480 450458 536
rect 450682 480 451654 536
rect 451878 480 452850 536
rect 453074 480 454046 536
rect 454270 480 455242 536
rect 455466 480 456346 536
rect 456570 480 457542 536
rect 457766 480 458738 536
rect 458962 480 459934 536
rect 460158 480 461038 536
rect 461262 480 462234 536
rect 462458 480 463430 536
rect 463654 480 464626 536
rect 464850 480 465730 536
rect 465954 480 466926 536
rect 467150 480 468122 536
rect 468346 480 469318 536
rect 469542 480 470514 536
rect 470738 480 471618 536
rect 471842 480 472814 536
rect 473038 480 474010 536
rect 474234 480 475206 536
rect 475430 480 476310 536
rect 476534 480 477506 536
rect 477730 480 478702 536
rect 478926 480 479898 536
rect 480122 480 481094 536
rect 481318 480 482198 536
rect 482422 480 483394 536
rect 483618 480 484590 536
rect 484814 480 485786 536
rect 486010 480 486890 536
rect 487114 480 488086 536
rect 488310 480 489282 536
rect 489506 480 490478 536
rect 490702 480 491582 536
rect 491806 480 492778 536
rect 493002 480 493974 536
rect 494198 480 495170 536
rect 495394 480 496366 536
rect 496590 480 497470 536
rect 497694 480 498666 536
rect 498890 480 499862 536
rect 500086 480 501058 536
rect 501282 480 502162 536
rect 502386 480 503358 536
rect 503582 480 504554 536
rect 504778 480 505750 536
rect 505974 480 506946 536
rect 507170 480 508050 536
rect 508274 480 509246 536
rect 509470 480 510442 536
rect 510666 480 511638 536
rect 511862 480 512742 536
rect 512966 480 513938 536
rect 514162 480 515134 536
rect 515358 480 516330 536
rect 516554 480 517434 536
rect 517658 480 518630 536
rect 518854 480 519826 536
rect 520050 480 521022 536
rect 521246 480 522218 536
rect 522442 480 523322 536
rect 523546 480 524518 536
rect 524742 480 525714 536
rect 525938 480 526910 536
rect 527134 480 528014 536
rect 528238 480 529210 536
rect 529434 480 530406 536
rect 530630 480 531602 536
rect 531826 480 532798 536
rect 533022 480 533902 536
rect 534126 480 535098 536
rect 535322 480 536294 536
rect 536518 480 537490 536
rect 537714 480 538594 536
rect 538818 480 539790 536
rect 540014 480 540986 536
rect 541210 480 542182 536
rect 542406 480 543286 536
rect 543510 480 544482 536
rect 544706 480 545678 536
rect 545902 480 546874 536
rect 547098 480 548070 536
rect 548294 480 549174 536
rect 549398 480 550370 536
rect 550594 480 551566 536
rect 551790 480 552762 536
rect 552986 480 553866 536
rect 554090 480 555062 536
rect 555286 480 556258 536
rect 556482 480 557454 536
rect 557678 480 558650 536
rect 558874 480 559754 536
rect 559978 480 560950 536
rect 561174 480 562146 536
rect 562370 480 563342 536
rect 563566 480 564446 536
rect 564670 480 565642 536
rect 565866 480 566838 536
rect 567062 480 568034 536
rect 568258 480 569138 536
rect 569362 480 570334 536
rect 570558 480 571530 536
rect 571754 480 572726 536
rect 572950 480 573922 536
rect 574146 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577418 536
rect 577642 480 578614 536
rect 578838 480 579718 536
rect 579942 480 580914 536
rect 581138 480 582110 536
rect 582334 480 583306 536
<< metal3 >>
rect 583520 698036 584960 698276
rect -960 697628 480 697868
rect 583520 686476 584960 686716
rect -960 685252 480 685492
rect 583520 674916 584960 675156
rect -960 672876 480 673116
rect 583520 663356 584960 663596
rect -960 660500 480 660740
rect 583520 651796 584960 652036
rect -960 648124 480 648364
rect 583520 640236 584960 640476
rect -960 635884 480 636124
rect 583520 628812 584960 629052
rect -960 623508 480 623748
rect 583520 617252 584960 617492
rect -960 611132 480 611372
rect 583520 605692 584960 605932
rect -960 598756 480 598996
rect 583520 594132 584960 594372
rect -960 586380 480 586620
rect 583520 582572 584960 582812
rect -960 574140 480 574380
rect 583520 571012 584960 571252
rect -960 561764 480 562004
rect 583520 559452 584960 559692
rect -960 549388 480 549628
rect 583520 548028 584960 548268
rect -960 537012 480 537252
rect 583520 536468 584960 536708
rect -960 524636 480 524876
rect 583520 524908 584960 525148
rect 583520 513348 584960 513588
rect -960 512396 480 512636
rect 583520 501788 584960 502028
rect -960 500020 480 500260
rect 583520 490228 584960 490468
rect -960 487644 480 487884
rect 583520 478668 584960 478908
rect -960 475268 480 475508
rect 583520 467244 584960 467484
rect -960 462892 480 463132
rect 583520 455684 584960 455924
rect -960 450652 480 450892
rect 583520 444124 584960 444364
rect -960 438276 480 438516
rect 583520 432564 584960 432804
rect -960 425900 480 426140
rect 583520 421004 584960 421244
rect -960 413524 480 413764
rect 583520 409444 584960 409684
rect -960 401148 480 401388
rect 583520 397884 584960 398124
rect -960 388908 480 389148
rect 583520 386460 584960 386700
rect -960 376532 480 376772
rect 583520 374900 584960 375140
rect -960 364156 480 364396
rect 583520 363340 584960 363580
rect -960 351780 480 352020
rect 583520 351780 584960 352020
rect 583520 340220 584960 340460
rect -960 339404 480 339644
rect 583520 328660 584960 328900
rect -960 327028 480 327268
rect 583520 317236 584960 317476
rect -960 314788 480 315028
rect 583520 305676 584960 305916
rect -960 302412 480 302652
rect 583520 294116 584960 294356
rect -960 290036 480 290276
rect 583520 282556 584960 282796
rect -960 277660 480 277900
rect 583520 270996 584960 271236
rect -960 265284 480 265524
rect 583520 259436 584960 259676
rect -960 253044 480 253284
rect 583520 247876 584960 248116
rect -960 240668 480 240908
rect 583520 236452 584960 236692
rect -960 228292 480 228532
rect 583520 224892 584960 225132
rect -960 215916 480 216156
rect 583520 213332 584960 213572
rect -960 203540 480 203780
rect 583520 201772 584960 202012
rect -960 191300 480 191540
rect 583520 190212 584960 190452
rect -960 178924 480 179164
rect 583520 178652 584960 178892
rect 583520 167092 584960 167332
rect -960 166548 480 166788
rect 583520 155668 584960 155908
rect -960 154172 480 154412
rect 583520 144108 584960 144348
rect -960 141796 480 142036
rect 583520 132548 584960 132788
rect -960 129556 480 129796
rect 583520 120988 584960 121228
rect -960 117180 480 117420
rect 583520 109428 584960 109668
rect -960 104804 480 105044
rect 583520 97868 584960 98108
rect -960 92428 480 92668
rect 583520 86308 584960 86548
rect -960 80052 480 80292
rect 583520 74884 584960 75124
rect -960 67812 480 68052
rect 583520 63324 584960 63564
rect -960 55436 480 55676
rect 583520 51764 584960 52004
rect -960 43060 480 43300
rect 583520 40204 584960 40444
rect -960 30684 480 30924
rect 583520 28644 584960 28884
rect -960 18308 480 18548
rect 583520 17084 584960 17324
rect -960 6068 480 6308
rect 583520 5660 584960 5900
<< obsm3 >>
rect 480 698356 583520 701793
rect 480 697956 583440 698356
rect 480 697948 583520 697956
rect 560 697548 583520 697948
rect 480 686796 583520 697548
rect 480 686396 583440 686796
rect 480 685572 583520 686396
rect 560 685172 583520 685572
rect 480 675236 583520 685172
rect 480 674836 583440 675236
rect 480 673196 583520 674836
rect 560 672796 583520 673196
rect 480 663676 583520 672796
rect 480 663276 583440 663676
rect 480 660820 583520 663276
rect 560 660420 583520 660820
rect 480 652116 583520 660420
rect 480 651716 583440 652116
rect 480 648444 583520 651716
rect 560 648044 583520 648444
rect 480 640556 583520 648044
rect 480 640156 583440 640556
rect 480 636204 583520 640156
rect 560 635804 583520 636204
rect 480 629132 583520 635804
rect 480 628732 583440 629132
rect 480 623828 583520 628732
rect 560 623428 583520 623828
rect 480 617572 583520 623428
rect 480 617172 583440 617572
rect 480 611452 583520 617172
rect 560 611052 583520 611452
rect 480 606012 583520 611052
rect 480 605612 583440 606012
rect 480 599076 583520 605612
rect 560 598676 583520 599076
rect 480 594452 583520 598676
rect 480 594052 583440 594452
rect 480 586700 583520 594052
rect 560 586300 583520 586700
rect 480 582892 583520 586300
rect 480 582492 583440 582892
rect 480 574460 583520 582492
rect 560 574060 583520 574460
rect 480 571332 583520 574060
rect 480 570932 583440 571332
rect 480 562084 583520 570932
rect 560 561684 583520 562084
rect 480 559772 583520 561684
rect 480 559372 583440 559772
rect 480 549708 583520 559372
rect 560 549308 583520 549708
rect 480 548348 583520 549308
rect 480 547948 583440 548348
rect 480 537332 583520 547948
rect 560 536932 583520 537332
rect 480 536788 583520 536932
rect 480 536388 583440 536788
rect 480 525228 583520 536388
rect 480 524956 583440 525228
rect 560 524828 583440 524956
rect 560 524556 583520 524828
rect 480 513668 583520 524556
rect 480 513268 583440 513668
rect 480 512716 583520 513268
rect 560 512316 583520 512716
rect 480 502108 583520 512316
rect 480 501708 583440 502108
rect 480 500340 583520 501708
rect 560 499940 583520 500340
rect 480 490548 583520 499940
rect 480 490148 583440 490548
rect 480 487964 583520 490148
rect 560 487564 583520 487964
rect 480 478988 583520 487564
rect 480 478588 583440 478988
rect 480 475588 583520 478588
rect 560 475188 583520 475588
rect 480 467564 583520 475188
rect 480 467164 583440 467564
rect 480 463212 583520 467164
rect 560 462812 583520 463212
rect 480 456004 583520 462812
rect 480 455604 583440 456004
rect 480 450972 583520 455604
rect 560 450572 583520 450972
rect 480 444444 583520 450572
rect 480 444044 583440 444444
rect 480 438596 583520 444044
rect 560 438196 583520 438596
rect 480 432884 583520 438196
rect 480 432484 583440 432884
rect 480 426220 583520 432484
rect 560 425820 583520 426220
rect 480 421324 583520 425820
rect 480 420924 583440 421324
rect 480 413844 583520 420924
rect 560 413444 583520 413844
rect 480 409764 583520 413444
rect 480 409364 583440 409764
rect 480 401468 583520 409364
rect 560 401068 583520 401468
rect 480 398204 583520 401068
rect 480 397804 583440 398204
rect 480 389228 583520 397804
rect 560 388828 583520 389228
rect 480 386780 583520 388828
rect 480 386380 583440 386780
rect 480 376852 583520 386380
rect 560 376452 583520 376852
rect 480 375220 583520 376452
rect 480 374820 583440 375220
rect 480 364476 583520 374820
rect 560 364076 583520 364476
rect 480 363660 583520 364076
rect 480 363260 583440 363660
rect 480 352100 583520 363260
rect 560 351700 583440 352100
rect 480 340540 583520 351700
rect 480 340140 583440 340540
rect 480 339724 583520 340140
rect 560 339324 583520 339724
rect 480 328980 583520 339324
rect 480 328580 583440 328980
rect 480 327348 583520 328580
rect 560 326948 583520 327348
rect 480 317556 583520 326948
rect 480 317156 583440 317556
rect 480 315108 583520 317156
rect 560 314708 583520 315108
rect 480 305996 583520 314708
rect 480 305596 583440 305996
rect 480 302732 583520 305596
rect 560 302332 583520 302732
rect 480 294436 583520 302332
rect 480 294036 583440 294436
rect 480 290356 583520 294036
rect 560 289956 583520 290356
rect 480 282876 583520 289956
rect 480 282476 583440 282876
rect 480 277980 583520 282476
rect 560 277580 583520 277980
rect 480 271316 583520 277580
rect 480 270916 583440 271316
rect 480 265604 583520 270916
rect 560 265204 583520 265604
rect 480 259756 583520 265204
rect 480 259356 583440 259756
rect 480 253364 583520 259356
rect 560 252964 583520 253364
rect 480 248196 583520 252964
rect 480 247796 583440 248196
rect 480 240988 583520 247796
rect 560 240588 583520 240988
rect 480 236772 583520 240588
rect 480 236372 583440 236772
rect 480 228612 583520 236372
rect 560 228212 583520 228612
rect 480 225212 583520 228212
rect 480 224812 583440 225212
rect 480 216236 583520 224812
rect 560 215836 583520 216236
rect 480 213652 583520 215836
rect 480 213252 583440 213652
rect 480 203860 583520 213252
rect 560 203460 583520 203860
rect 480 202092 583520 203460
rect 480 201692 583440 202092
rect 480 191620 583520 201692
rect 560 191220 583520 191620
rect 480 190532 583520 191220
rect 480 190132 583440 190532
rect 480 179244 583520 190132
rect 560 178972 583520 179244
rect 560 178844 583440 178972
rect 480 178572 583440 178844
rect 480 167412 583520 178572
rect 480 167012 583440 167412
rect 480 166868 583520 167012
rect 560 166468 583520 166868
rect 480 155988 583520 166468
rect 480 155588 583440 155988
rect 480 154492 583520 155588
rect 560 154092 583520 154492
rect 480 144428 583520 154092
rect 480 144028 583440 144428
rect 480 142116 583520 144028
rect 560 141716 583520 142116
rect 480 132868 583520 141716
rect 480 132468 583440 132868
rect 480 129876 583520 132468
rect 560 129476 583520 129876
rect 480 121308 583520 129476
rect 480 120908 583440 121308
rect 480 117500 583520 120908
rect 560 117100 583520 117500
rect 480 109748 583520 117100
rect 480 109348 583440 109748
rect 480 105124 583520 109348
rect 560 104724 583520 105124
rect 480 98188 583520 104724
rect 480 97788 583440 98188
rect 480 92748 583520 97788
rect 560 92348 583520 92748
rect 480 86628 583520 92348
rect 480 86228 583440 86628
rect 480 80372 583520 86228
rect 560 79972 583520 80372
rect 480 75204 583520 79972
rect 480 74804 583440 75204
rect 480 68132 583520 74804
rect 560 67732 583520 68132
rect 480 63644 583520 67732
rect 480 63244 583440 63644
rect 480 55756 583520 63244
rect 560 55356 583520 55756
rect 480 52084 583520 55356
rect 480 51684 583440 52084
rect 480 43380 583520 51684
rect 560 42980 583520 43380
rect 480 40524 583520 42980
rect 480 40124 583440 40524
rect 480 31004 583520 40124
rect 560 30604 583520 31004
rect 480 28964 583520 30604
rect 480 28564 583440 28964
rect 480 18628 583520 28564
rect 560 18228 583520 18628
rect 480 17404 583520 18228
rect 480 17004 583440 17404
rect 480 6388 583520 17004
rect 560 5988 583520 6388
rect 480 5980 583520 5988
rect 480 5580 583440 5980
rect 480 2143 583520 5580
<< metal4 >>
rect -8576 -7504 -7976 711440
rect -7636 -6564 -7036 710500
rect -6696 -5624 -6096 709560
rect -5756 -4684 -5156 708620
rect -4816 -3744 -4216 707680
rect -3876 -2804 -3276 706740
rect -2936 -1864 -2336 705800
rect -1996 -924 -1396 704860
rect 1804 -1864 2404 705800
rect 5404 -3744 6004 707680
rect 9004 -5624 9604 709560
rect 12604 -7504 13204 711440
rect 19804 -1864 20404 705800
rect 23404 -3744 24004 707680
rect 27004 -5624 27604 709560
rect 30604 -7504 31204 711440
rect 37804 -1864 38404 705800
rect 41404 -3744 42004 707680
rect 45004 -5624 45604 709560
rect 48604 -7504 49204 711440
rect 55804 -1864 56404 705800
rect 59404 -3744 60004 707680
rect 63004 -5624 63604 709560
rect 66604 -7504 67204 711440
rect 73804 -1864 74404 705800
rect 77404 -3744 78004 707680
rect 81004 -5624 81604 709560
rect 84604 -7504 85204 711440
rect 91804 -1864 92404 705800
rect 95404 -3744 96004 707680
rect 99004 -5624 99604 709560
rect 102604 -7504 103204 711440
rect 109804 -1864 110404 705800
rect 113404 -3744 114004 707680
rect 117004 -5624 117604 709560
rect 120604 -7504 121204 711440
rect 127804 -1864 128404 705800
rect 131404 -3744 132004 707680
rect 135004 -5624 135604 709560
rect 138604 -7504 139204 711440
rect 145804 -1864 146404 705800
rect 149404 -3744 150004 707680
rect 153004 -5624 153604 709560
rect 156604 -7504 157204 711440
rect 163804 -1864 164404 705800
rect 167404 -3744 168004 707680
rect 171004 -5624 171604 709560
rect 174604 -7504 175204 711440
rect 181804 -1864 182404 705800
rect 185404 -3744 186004 707680
rect 189004 -5624 189604 709560
rect 192604 -7504 193204 711440
rect 199804 -1864 200404 705800
rect 203404 -3744 204004 707680
rect 207004 -5624 207604 709560
rect 210604 -7504 211204 711440
rect 217804 -1864 218404 705800
rect 221404 -3744 222004 707680
rect 225004 -5624 225604 709560
rect 228604 -7504 229204 711440
rect 235804 459952 236404 705800
rect 239404 460000 240004 707680
rect 243004 460000 243604 709560
rect 246604 460000 247204 711440
rect 253804 459952 254404 705800
rect 257404 460000 258004 707680
rect 261004 460000 261604 709560
rect 264604 460000 265204 711440
rect 271804 459952 272404 705800
rect 275404 460000 276004 707680
rect 279004 460000 279604 709560
rect 282604 460000 283204 711440
rect 289804 459952 290404 705800
rect 293404 460000 294004 707680
rect 297004 460000 297604 709560
rect 300604 460000 301204 711440
rect 307804 459952 308404 705800
rect 311404 460000 312004 707680
rect 315004 460000 315604 709560
rect 318604 460000 319204 711440
rect 325804 459952 326404 705800
rect 329404 460000 330004 707680
rect 333004 460000 333604 709560
rect 336604 460000 337204 711440
rect 343804 459952 344404 705800
rect 347404 460000 348004 707680
rect 351004 460000 351604 709560
rect 354604 460000 355204 711440
rect 235804 -1864 236404 336048
rect 239404 -3744 240004 336000
rect 243004 -5624 243604 336000
rect 246604 -7504 247204 336000
rect 253804 -1864 254404 336048
rect 257404 -3744 258004 336000
rect 261004 -5624 261604 336000
rect 264604 -7504 265204 336000
rect 271804 -1864 272404 336048
rect 275404 -3744 276004 336000
rect 279004 -5624 279604 336000
rect 282604 -7504 283204 336000
rect 289804 -1864 290404 336048
rect 293404 -3744 294004 336000
rect 297004 -5624 297604 336000
rect 300604 -7504 301204 336000
rect 307804 -1864 308404 336048
rect 311404 -3744 312004 336000
rect 315004 -5624 315604 336000
rect 318604 -7504 319204 336000
rect 325804 -1864 326404 336048
rect 329404 -3744 330004 336000
rect 333004 -5624 333604 336000
rect 336604 -7504 337204 336000
rect 343804 -1864 344404 336048
rect 347404 -3744 348004 336000
rect 351004 -5624 351604 336000
rect 354604 -7504 355204 336000
rect 361804 -1864 362404 705800
rect 365404 -3744 366004 707680
rect 369004 -5624 369604 709560
rect 372604 -7504 373204 711440
rect 379804 -1864 380404 705800
rect 383404 -3744 384004 707680
rect 387004 -5624 387604 709560
rect 390604 -7504 391204 711440
rect 397804 -1864 398404 705800
rect 401404 -3744 402004 707680
rect 405004 -5624 405604 709560
rect 408604 -7504 409204 711440
rect 415804 -1864 416404 705800
rect 419404 -3744 420004 707680
rect 423004 -5624 423604 709560
rect 426604 -7504 427204 711440
rect 433804 -1864 434404 705800
rect 437404 -3744 438004 707680
rect 441004 -5624 441604 709560
rect 444604 -7504 445204 711440
rect 451804 -1864 452404 705800
rect 455404 -3744 456004 707680
rect 459004 -5624 459604 709560
rect 462604 -7504 463204 711440
rect 469804 -1864 470404 705800
rect 473404 -3744 474004 707680
rect 477004 -5624 477604 709560
rect 480604 -7504 481204 711440
rect 487804 -1864 488404 705800
rect 491404 -3744 492004 707680
rect 495004 -5624 495604 709560
rect 498604 -7504 499204 711440
rect 505804 -1864 506404 705800
rect 509404 -3744 510004 707680
rect 513004 -5624 513604 709560
rect 516604 -7504 517204 711440
rect 523804 -1864 524404 705800
rect 527404 -3744 528004 707680
rect 531004 -5624 531604 709560
rect 534604 -7504 535204 711440
rect 541804 -1864 542404 705800
rect 545404 -3744 546004 707680
rect 549004 -5624 549604 709560
rect 552604 -7504 553204 711440
rect 559804 -1864 560404 705800
rect 563404 -3744 564004 707680
rect 567004 -5624 567604 709560
rect 570604 -7504 571204 711440
rect 577804 -1864 578404 705800
rect 581404 -3744 582004 707680
rect 585320 -924 585920 704860
rect 586260 -1864 586860 705800
rect 587200 -2804 587800 706740
rect 588140 -3744 588740 707680
rect 589080 -4684 589680 708620
rect 590020 -5624 590620 709560
rect 590960 -6564 591560 710500
rect 591900 -7504 592500 711440
<< obsm4 >>
rect 237235 336128 361724 457469
rect 237235 336080 253724 336128
rect 237235 6835 239324 336080
rect 240084 6835 242924 336080
rect 243684 6835 246524 336080
rect 247284 6835 253724 336080
rect 254484 336080 271724 336128
rect 254484 6835 257324 336080
rect 258084 6835 260924 336080
rect 261684 6835 264524 336080
rect 265284 6835 271724 336080
rect 272484 336080 289724 336128
rect 272484 6835 275324 336080
rect 276084 6835 278924 336080
rect 279684 6835 282524 336080
rect 283284 6835 289724 336080
rect 290484 336080 307724 336128
rect 290484 6835 293324 336080
rect 294084 6835 296924 336080
rect 297684 6835 300524 336080
rect 301284 6835 307724 336080
rect 308484 336080 325724 336128
rect 308484 6835 311324 336080
rect 312084 6835 314924 336080
rect 315684 6835 318524 336080
rect 319284 6835 325724 336080
rect 326484 336080 343724 336128
rect 326484 6835 329324 336080
rect 330084 6835 332924 336080
rect 333684 6835 336524 336080
rect 337284 6835 343724 336080
rect 344484 336080 361724 336128
rect 344484 6835 347324 336080
rect 348084 6835 350924 336080
rect 351684 6835 354524 336080
rect 355284 6835 361724 336080
rect 362484 6835 365324 457469
rect 366084 6835 368924 457469
rect 369684 6835 372524 457469
rect 373284 6835 379724 457469
rect 380484 6835 383324 457469
rect 384084 6835 386924 457469
rect 387684 6835 390524 457469
rect 391284 6835 397724 457469
rect 398484 6835 401324 457469
rect 402084 6835 404924 457469
rect 405684 6835 408524 457469
rect 409284 6835 415724 457469
rect 416484 6835 419324 457469
rect 420084 6835 422924 457469
rect 423684 6835 426524 457469
rect 427284 6835 433724 457469
rect 434484 6835 437324 457469
rect 438084 6835 440924 457469
rect 441684 6835 444524 457469
rect 445284 6835 451724 457469
rect 452484 6835 455324 457469
rect 456084 6835 458924 457469
rect 459684 6835 462524 457469
rect 463284 6835 469724 457469
rect 470484 6835 473324 457469
rect 474084 6835 476924 457469
rect 477684 6835 480524 457469
rect 481284 6835 487724 457469
rect 488484 6835 491324 457469
rect 492084 6835 494924 457469
rect 495684 6835 498524 457469
rect 499284 6835 505724 457469
rect 506484 6835 509324 457469
rect 510084 6835 512924 457469
rect 513684 6835 516524 457469
rect 517284 6835 523724 457469
rect 524484 6835 527324 457469
rect 528084 6835 530924 457469
rect 531684 6835 534524 457469
rect 535284 6835 541724 457469
rect 542484 6835 545324 457469
rect 546084 6835 548924 457469
rect 549684 6835 552524 457469
rect 553284 6835 559724 457469
rect 560484 6835 563324 457469
rect 564084 6835 566924 457469
rect 567684 6835 570524 457469
rect 571284 6835 577724 457469
rect 578484 6835 580362 457469
<< metal5 >>
rect -8576 710840 592500 711440
rect -7636 709900 591560 710500
rect -6696 708960 590620 709560
rect -5756 708020 589680 708620
rect -4816 707080 588740 707680
rect -3876 706140 587800 706740
rect -2936 705200 586860 705800
rect -1996 704260 585920 704860
rect -8576 697676 592500 698276
rect -6696 694076 590620 694676
rect -4816 690476 588740 691076
rect -2936 686828 586860 687428
rect -8576 679676 592500 680276
rect -6696 676076 590620 676676
rect -4816 672476 588740 673076
rect -2936 668828 586860 669428
rect -8576 661676 592500 662276
rect -6696 658076 590620 658676
rect -4816 654476 588740 655076
rect -2936 650828 586860 651428
rect -8576 643676 592500 644276
rect -6696 640076 590620 640676
rect -4816 636476 588740 637076
rect -2936 632828 586860 633428
rect -8576 625676 592500 626276
rect -6696 622076 590620 622676
rect -4816 618476 588740 619076
rect -2936 614828 586860 615428
rect -8576 607676 592500 608276
rect -6696 604076 590620 604676
rect -4816 600476 588740 601076
rect -2936 596828 586860 597428
rect -8576 589676 592500 590276
rect -6696 586076 590620 586676
rect -4816 582476 588740 583076
rect -2936 578828 586860 579428
rect -8576 571676 592500 572276
rect -6696 568076 590620 568676
rect -4816 564476 588740 565076
rect -2936 560828 586860 561428
rect -8576 553676 592500 554276
rect -6696 550076 590620 550676
rect -4816 546476 588740 547076
rect -2936 542828 586860 543428
rect -8576 535676 592500 536276
rect -6696 532076 590620 532676
rect -4816 528476 588740 529076
rect -2936 524828 586860 525428
rect -8576 517676 592500 518276
rect -6696 514076 590620 514676
rect -4816 510476 588740 511076
rect -2936 506828 586860 507428
rect -8576 499676 592500 500276
rect -6696 496076 590620 496676
rect -4816 492476 588740 493076
rect -2936 488828 586860 489428
rect -8576 481676 592500 482276
rect -6696 478076 590620 478676
rect -4816 474476 588740 475076
rect -2936 470828 586860 471428
rect -8576 463676 592500 464276
rect -6696 460076 590620 460676
rect -4816 456476 588740 457076
rect -2936 452828 586860 453428
rect -8576 445676 592500 446276
rect -6696 442076 590620 442676
rect -4816 438476 588740 439076
rect -2936 434828 586860 435428
rect -8576 427676 592500 428276
rect -6696 424076 590620 424676
rect -4816 420476 588740 421076
rect -2936 416828 586860 417428
rect -8576 409676 592500 410276
rect -6696 406076 590620 406676
rect -4816 402476 588740 403076
rect -2936 398828 586860 399428
rect -8576 391676 592500 392276
rect -6696 388076 590620 388676
rect -4816 384476 588740 385076
rect -2936 380828 586860 381428
rect -8576 373676 592500 374276
rect -6696 370076 590620 370676
rect -4816 366476 588740 367076
rect -2936 362828 586860 363428
rect -8576 355676 592500 356276
rect -6696 352076 590620 352676
rect -4816 348476 588740 349076
rect -2936 344828 586860 345428
rect -8576 337676 592500 338276
rect -6696 334076 590620 334676
rect -4816 330476 588740 331076
rect -2936 326828 586860 327428
rect -8576 319676 592500 320276
rect -6696 316076 590620 316676
rect -4816 312476 588740 313076
rect -2936 308828 586860 309428
rect -8576 301676 592500 302276
rect -6696 298076 590620 298676
rect -4816 294476 588740 295076
rect -2936 290828 586860 291428
rect -8576 283676 592500 284276
rect -6696 280076 590620 280676
rect -4816 276476 588740 277076
rect -2936 272828 586860 273428
rect -8576 265676 592500 266276
rect -6696 262076 590620 262676
rect -4816 258476 588740 259076
rect -2936 254828 586860 255428
rect -8576 247676 592500 248276
rect -6696 244076 590620 244676
rect -4816 240476 588740 241076
rect -2936 236828 586860 237428
rect -8576 229676 592500 230276
rect -6696 226076 590620 226676
rect -4816 222476 588740 223076
rect -2936 218828 586860 219428
rect -8576 211676 592500 212276
rect -6696 208076 590620 208676
rect -4816 204476 588740 205076
rect -2936 200828 586860 201428
rect -8576 193676 592500 194276
rect -6696 190076 590620 190676
rect -4816 186476 588740 187076
rect -2936 182828 586860 183428
rect -8576 175676 592500 176276
rect -6696 172076 590620 172676
rect -4816 168476 588740 169076
rect -2936 164828 586860 165428
rect -8576 157676 592500 158276
rect -6696 154076 590620 154676
rect -4816 150476 588740 151076
rect -2936 146828 586860 147428
rect -8576 139676 592500 140276
rect -6696 136076 590620 136676
rect -4816 132476 588740 133076
rect -2936 128828 586860 129428
rect -8576 121676 592500 122276
rect -6696 118076 590620 118676
rect -4816 114476 588740 115076
rect -2936 110828 586860 111428
rect -8576 103676 592500 104276
rect -6696 100076 590620 100676
rect -4816 96476 588740 97076
rect -2936 92828 586860 93428
rect -8576 85676 592500 86276
rect -6696 82076 590620 82676
rect -4816 78476 588740 79076
rect -2936 74828 586860 75428
rect -8576 67676 592500 68276
rect -6696 64076 590620 64676
rect -4816 60476 588740 61076
rect -2936 56828 586860 57428
rect -8576 49676 592500 50276
rect -6696 46076 590620 46676
rect -4816 42476 588740 43076
rect -2936 38828 586860 39428
rect -8576 31676 592500 32276
rect -6696 28076 590620 28676
rect -4816 24476 588740 25076
rect -2936 20828 586860 21428
rect -8576 13676 592500 14276
rect -6696 10076 590620 10676
rect -4816 6476 588740 7076
rect -2936 2828 586860 3428
rect -1996 -924 585920 -324
rect -2936 -1864 586860 -1264
rect -3876 -2804 587800 -2204
rect -4816 -3744 588740 -3144
rect -5756 -4684 589680 -4084
rect -6696 -5624 590620 -5024
rect -7636 -6564 591560 -5964
rect -8576 -7504 592500 -6904
<< obsm5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect 0 698596 584000 703940
rect -7636 698276 -7036 698278
rect 590960 698276 591560 698278
rect -7636 697674 -7036 697676
rect 590960 697674 591560 697676
rect 0 694996 584000 697356
rect -5756 694676 -5156 694678
rect 589080 694676 589680 694678
rect -5756 694074 -5156 694076
rect 589080 694074 589680 694076
rect 0 691396 584000 693756
rect -3876 691076 -3276 691078
rect 587200 691076 587800 691078
rect -3876 690474 -3276 690476
rect 587200 690474 587800 690476
rect 0 687748 584000 690156
rect -1996 687428 -1396 687430
rect 585320 687428 585920 687430
rect -1996 686826 -1396 686828
rect 585320 686826 585920 686828
rect 0 680596 584000 686508
rect -8576 680276 -7976 680278
rect 591900 680276 592500 680278
rect -8576 679674 -7976 679676
rect 591900 679674 592500 679676
rect 0 676996 584000 679356
rect -6696 676676 -6096 676678
rect 590020 676676 590620 676678
rect -6696 676074 -6096 676076
rect 590020 676074 590620 676076
rect 0 673396 584000 675756
rect -4816 673076 -4216 673078
rect 588140 673076 588740 673078
rect -4816 672474 -4216 672476
rect 588140 672474 588740 672476
rect 0 669748 584000 672156
rect -2936 669428 -2336 669430
rect 586260 669428 586860 669430
rect -2936 668826 -2336 668828
rect 586260 668826 586860 668828
rect 0 662596 584000 668508
rect -7636 662276 -7036 662278
rect 590960 662276 591560 662278
rect -7636 661674 -7036 661676
rect 590960 661674 591560 661676
rect 0 658996 584000 661356
rect -5756 658676 -5156 658678
rect 589080 658676 589680 658678
rect -5756 658074 -5156 658076
rect 589080 658074 589680 658076
rect 0 655396 584000 657756
rect -3876 655076 -3276 655078
rect 587200 655076 587800 655078
rect -3876 654474 -3276 654476
rect 587200 654474 587800 654476
rect 0 651748 584000 654156
rect -1996 651428 -1396 651430
rect 585320 651428 585920 651430
rect -1996 650826 -1396 650828
rect 585320 650826 585920 650828
rect 0 644596 584000 650508
rect -8576 644276 -7976 644278
rect 591900 644276 592500 644278
rect -8576 643674 -7976 643676
rect 591900 643674 592500 643676
rect 0 640996 584000 643356
rect -6696 640676 -6096 640678
rect 590020 640676 590620 640678
rect -6696 640074 -6096 640076
rect 590020 640074 590620 640076
rect 0 637396 584000 639756
rect -4816 637076 -4216 637078
rect 588140 637076 588740 637078
rect -4816 636474 -4216 636476
rect 588140 636474 588740 636476
rect 0 633748 584000 636156
rect -2936 633428 -2336 633430
rect 586260 633428 586860 633430
rect -2936 632826 -2336 632828
rect 586260 632826 586860 632828
rect 0 626596 584000 632508
rect -7636 626276 -7036 626278
rect 590960 626276 591560 626278
rect -7636 625674 -7036 625676
rect 590960 625674 591560 625676
rect 0 622996 584000 625356
rect -5756 622676 -5156 622678
rect 589080 622676 589680 622678
rect -5756 622074 -5156 622076
rect 589080 622074 589680 622076
rect 0 619396 584000 621756
rect -3876 619076 -3276 619078
rect 587200 619076 587800 619078
rect -3876 618474 -3276 618476
rect 587200 618474 587800 618476
rect 0 615748 584000 618156
rect -1996 615428 -1396 615430
rect 585320 615428 585920 615430
rect -1996 614826 -1396 614828
rect 585320 614826 585920 614828
rect 0 608596 584000 614508
rect -8576 608276 -7976 608278
rect 591900 608276 592500 608278
rect -8576 607674 -7976 607676
rect 591900 607674 592500 607676
rect 0 604996 584000 607356
rect -6696 604676 -6096 604678
rect 590020 604676 590620 604678
rect -6696 604074 -6096 604076
rect 590020 604074 590620 604076
rect 0 601396 584000 603756
rect -4816 601076 -4216 601078
rect 588140 601076 588740 601078
rect -4816 600474 -4216 600476
rect 588140 600474 588740 600476
rect 0 597748 584000 600156
rect -2936 597428 -2336 597430
rect 586260 597428 586860 597430
rect -2936 596826 -2336 596828
rect 586260 596826 586860 596828
rect 0 590596 584000 596508
rect -7636 590276 -7036 590278
rect 590960 590276 591560 590278
rect -7636 589674 -7036 589676
rect 590960 589674 591560 589676
rect 0 586996 584000 589356
rect -5756 586676 -5156 586678
rect 589080 586676 589680 586678
rect -5756 586074 -5156 586076
rect 589080 586074 589680 586076
rect 0 583396 584000 585756
rect -3876 583076 -3276 583078
rect 587200 583076 587800 583078
rect -3876 582474 -3276 582476
rect 587200 582474 587800 582476
rect 0 579748 584000 582156
rect -1996 579428 -1396 579430
rect 585320 579428 585920 579430
rect -1996 578826 -1396 578828
rect 585320 578826 585920 578828
rect 0 572596 584000 578508
rect -8576 572276 -7976 572278
rect 591900 572276 592500 572278
rect -8576 571674 -7976 571676
rect 591900 571674 592500 571676
rect 0 568996 584000 571356
rect -6696 568676 -6096 568678
rect 590020 568676 590620 568678
rect -6696 568074 -6096 568076
rect 590020 568074 590620 568076
rect 0 565396 584000 567756
rect -4816 565076 -4216 565078
rect 588140 565076 588740 565078
rect -4816 564474 -4216 564476
rect 588140 564474 588740 564476
rect 0 561748 584000 564156
rect -2936 561428 -2336 561430
rect 586260 561428 586860 561430
rect -2936 560826 -2336 560828
rect 586260 560826 586860 560828
rect 0 554596 584000 560508
rect -7636 554276 -7036 554278
rect 590960 554276 591560 554278
rect -7636 553674 -7036 553676
rect 590960 553674 591560 553676
rect 0 550996 584000 553356
rect -5756 550676 -5156 550678
rect 589080 550676 589680 550678
rect -5756 550074 -5156 550076
rect 589080 550074 589680 550076
rect 0 547396 584000 549756
rect -3876 547076 -3276 547078
rect 587200 547076 587800 547078
rect -3876 546474 -3276 546476
rect 587200 546474 587800 546476
rect 0 543748 584000 546156
rect -1996 543428 -1396 543430
rect 585320 543428 585920 543430
rect -1996 542826 -1396 542828
rect 585320 542826 585920 542828
rect 0 536596 584000 542508
rect -8576 536276 -7976 536278
rect 591900 536276 592500 536278
rect -8576 535674 -7976 535676
rect 591900 535674 592500 535676
rect 0 532996 584000 535356
rect -6696 532676 -6096 532678
rect 590020 532676 590620 532678
rect -6696 532074 -6096 532076
rect 590020 532074 590620 532076
rect 0 529396 584000 531756
rect -4816 529076 -4216 529078
rect 588140 529076 588740 529078
rect -4816 528474 -4216 528476
rect 588140 528474 588740 528476
rect 0 525748 584000 528156
rect -2936 525428 -2336 525430
rect 586260 525428 586860 525430
rect -2936 524826 -2336 524828
rect 586260 524826 586860 524828
rect 0 518596 584000 524508
rect -7636 518276 -7036 518278
rect 590960 518276 591560 518278
rect -7636 517674 -7036 517676
rect 590960 517674 591560 517676
rect 0 514996 584000 517356
rect -5756 514676 -5156 514678
rect 589080 514676 589680 514678
rect -5756 514074 -5156 514076
rect 589080 514074 589680 514076
rect 0 511396 584000 513756
rect -3876 511076 -3276 511078
rect 587200 511076 587800 511078
rect -3876 510474 -3276 510476
rect 587200 510474 587800 510476
rect 0 507748 584000 510156
rect -1996 507428 -1396 507430
rect 585320 507428 585920 507430
rect -1996 506826 -1396 506828
rect 585320 506826 585920 506828
rect 0 500596 584000 506508
rect -8576 500276 -7976 500278
rect 591900 500276 592500 500278
rect -8576 499674 -7976 499676
rect 591900 499674 592500 499676
rect 0 496996 584000 499356
rect -6696 496676 -6096 496678
rect 590020 496676 590620 496678
rect -6696 496074 -6096 496076
rect 590020 496074 590620 496076
rect 0 493396 584000 495756
rect -4816 493076 -4216 493078
rect 588140 493076 588740 493078
rect -4816 492474 -4216 492476
rect 588140 492474 588740 492476
rect 0 489748 584000 492156
rect -2936 489428 -2336 489430
rect 586260 489428 586860 489430
rect -2936 488826 -2336 488828
rect 586260 488826 586860 488828
rect 0 482596 584000 488508
rect -7636 482276 -7036 482278
rect 590960 482276 591560 482278
rect -7636 481674 -7036 481676
rect 590960 481674 591560 481676
rect 0 478996 584000 481356
rect -5756 478676 -5156 478678
rect 589080 478676 589680 478678
rect -5756 478074 -5156 478076
rect 589080 478074 589680 478076
rect 0 475396 584000 477756
rect -3876 475076 -3276 475078
rect 587200 475076 587800 475078
rect -3876 474474 -3276 474476
rect 587200 474474 587800 474476
rect 0 471748 584000 474156
rect -1996 471428 -1396 471430
rect 585320 471428 585920 471430
rect -1996 470826 -1396 470828
rect 585320 470826 585920 470828
rect 0 464596 584000 470508
rect -8576 464276 -7976 464278
rect 591900 464276 592500 464278
rect -8576 463674 -7976 463676
rect 591900 463674 592500 463676
rect 0 460996 584000 463356
rect -6696 460676 -6096 460678
rect 590020 460676 590620 460678
rect -6696 460074 -6096 460076
rect 590020 460074 590620 460076
rect 0 457396 584000 459756
rect -4816 457076 -4216 457078
rect 588140 457076 588740 457078
rect -4816 456474 -4216 456476
rect 588140 456474 588740 456476
rect 0 453748 584000 456156
rect -2936 453428 -2336 453430
rect 586260 453428 586860 453430
rect -2936 452826 -2336 452828
rect 586260 452826 586860 452828
rect 0 446596 584000 452508
rect -7636 446276 -7036 446278
rect 590960 446276 591560 446278
rect -7636 445674 -7036 445676
rect 590960 445674 591560 445676
rect 0 442996 584000 445356
rect -5756 442676 -5156 442678
rect 589080 442676 589680 442678
rect -5756 442074 -5156 442076
rect 589080 442074 589680 442076
rect 0 439396 584000 441756
rect -3876 439076 -3276 439078
rect 587200 439076 587800 439078
rect -3876 438474 -3276 438476
rect 587200 438474 587800 438476
rect 0 435748 584000 438156
rect -1996 435428 -1396 435430
rect 585320 435428 585920 435430
rect -1996 434826 -1396 434828
rect 585320 434826 585920 434828
rect 0 428596 584000 434508
rect -8576 428276 -7976 428278
rect 591900 428276 592500 428278
rect -8576 427674 -7976 427676
rect 591900 427674 592500 427676
rect 0 424996 584000 427356
rect -6696 424676 -6096 424678
rect 590020 424676 590620 424678
rect -6696 424074 -6096 424076
rect 590020 424074 590620 424076
rect 0 421396 584000 423756
rect -4816 421076 -4216 421078
rect 588140 421076 588740 421078
rect -4816 420474 -4216 420476
rect 588140 420474 588740 420476
rect 0 417748 584000 420156
rect -2936 417428 -2336 417430
rect 586260 417428 586860 417430
rect -2936 416826 -2336 416828
rect 586260 416826 586860 416828
rect 0 410596 584000 416508
rect -7636 410276 -7036 410278
rect 590960 410276 591560 410278
rect -7636 409674 -7036 409676
rect 590960 409674 591560 409676
rect 0 406996 584000 409356
rect -5756 406676 -5156 406678
rect 589080 406676 589680 406678
rect -5756 406074 -5156 406076
rect 589080 406074 589680 406076
rect 0 403396 584000 405756
rect -3876 403076 -3276 403078
rect 587200 403076 587800 403078
rect -3876 402474 -3276 402476
rect 587200 402474 587800 402476
rect 0 399748 584000 402156
rect -1996 399428 -1396 399430
rect 585320 399428 585920 399430
rect -1996 398826 -1396 398828
rect 585320 398826 585920 398828
rect 0 392596 584000 398508
rect -8576 392276 -7976 392278
rect 591900 392276 592500 392278
rect -8576 391674 -7976 391676
rect 591900 391674 592500 391676
rect 0 388996 584000 391356
rect -6696 388676 -6096 388678
rect 590020 388676 590620 388678
rect -6696 388074 -6096 388076
rect 590020 388074 590620 388076
rect 0 385396 584000 387756
rect -4816 385076 -4216 385078
rect 588140 385076 588740 385078
rect -4816 384474 -4216 384476
rect 588140 384474 588740 384476
rect 0 381748 584000 384156
rect -2936 381428 -2336 381430
rect 586260 381428 586860 381430
rect -2936 380826 -2336 380828
rect 586260 380826 586860 380828
rect 0 374596 584000 380508
rect -7636 374276 -7036 374278
rect 590960 374276 591560 374278
rect -7636 373674 -7036 373676
rect 590960 373674 591560 373676
rect 0 370996 584000 373356
rect -5756 370676 -5156 370678
rect 589080 370676 589680 370678
rect -5756 370074 -5156 370076
rect 589080 370074 589680 370076
rect 0 367396 584000 369756
rect -3876 367076 -3276 367078
rect 587200 367076 587800 367078
rect -3876 366474 -3276 366476
rect 587200 366474 587800 366476
rect 0 363748 584000 366156
rect -1996 363428 -1396 363430
rect 585320 363428 585920 363430
rect -1996 362826 -1396 362828
rect 585320 362826 585920 362828
rect 0 356596 584000 362508
rect -8576 356276 -7976 356278
rect 591900 356276 592500 356278
rect -8576 355674 -7976 355676
rect 591900 355674 592500 355676
rect 0 352996 584000 355356
rect -6696 352676 -6096 352678
rect 590020 352676 590620 352678
rect -6696 352074 -6096 352076
rect 590020 352074 590620 352076
rect 0 349396 584000 351756
rect -4816 349076 -4216 349078
rect 588140 349076 588740 349078
rect -4816 348474 -4216 348476
rect 588140 348474 588740 348476
rect 0 345748 584000 348156
rect -2936 345428 -2336 345430
rect 586260 345428 586860 345430
rect -2936 344826 -2336 344828
rect 586260 344826 586860 344828
rect 0 338596 584000 344508
rect -7636 338276 -7036 338278
rect 590960 338276 591560 338278
rect -7636 337674 -7036 337676
rect 590960 337674 591560 337676
rect 0 334996 584000 337356
rect -5756 334676 -5156 334678
rect 589080 334676 589680 334678
rect -5756 334074 -5156 334076
rect 589080 334074 589680 334076
rect 0 331396 584000 333756
rect -3876 331076 -3276 331078
rect 587200 331076 587800 331078
rect -3876 330474 -3276 330476
rect 587200 330474 587800 330476
rect 0 327748 584000 330156
rect -1996 327428 -1396 327430
rect 585320 327428 585920 327430
rect -1996 326826 -1396 326828
rect 585320 326826 585920 326828
rect 0 320596 584000 326508
rect -8576 320276 -7976 320278
rect 591900 320276 592500 320278
rect -8576 319674 -7976 319676
rect 591900 319674 592500 319676
rect 0 316996 584000 319356
rect -6696 316676 -6096 316678
rect 590020 316676 590620 316678
rect -6696 316074 -6096 316076
rect 590020 316074 590620 316076
rect 0 313396 584000 315756
rect -4816 313076 -4216 313078
rect 588140 313076 588740 313078
rect -4816 312474 -4216 312476
rect 588140 312474 588740 312476
rect 0 309748 584000 312156
rect -2936 309428 -2336 309430
rect 586260 309428 586860 309430
rect -2936 308826 -2336 308828
rect 586260 308826 586860 308828
rect 0 302596 584000 308508
rect -7636 302276 -7036 302278
rect 590960 302276 591560 302278
rect -7636 301674 -7036 301676
rect 590960 301674 591560 301676
rect 0 298996 584000 301356
rect -5756 298676 -5156 298678
rect 589080 298676 589680 298678
rect -5756 298074 -5156 298076
rect 589080 298074 589680 298076
rect 0 295396 584000 297756
rect -3876 295076 -3276 295078
rect 587200 295076 587800 295078
rect -3876 294474 -3276 294476
rect 587200 294474 587800 294476
rect 0 291748 584000 294156
rect -1996 291428 -1396 291430
rect 585320 291428 585920 291430
rect -1996 290826 -1396 290828
rect 585320 290826 585920 290828
rect 0 284596 584000 290508
rect -8576 284276 -7976 284278
rect 591900 284276 592500 284278
rect -8576 283674 -7976 283676
rect 591900 283674 592500 283676
rect 0 280996 584000 283356
rect -6696 280676 -6096 280678
rect 590020 280676 590620 280678
rect -6696 280074 -6096 280076
rect 590020 280074 590620 280076
rect 0 277396 584000 279756
rect -4816 277076 -4216 277078
rect 588140 277076 588740 277078
rect -4816 276474 -4216 276476
rect 588140 276474 588740 276476
rect 0 273748 584000 276156
rect -2936 273428 -2336 273430
rect 586260 273428 586860 273430
rect -2936 272826 -2336 272828
rect 586260 272826 586860 272828
rect 0 266596 584000 272508
rect -7636 266276 -7036 266278
rect 590960 266276 591560 266278
rect -7636 265674 -7036 265676
rect 590960 265674 591560 265676
rect 0 262996 584000 265356
rect -5756 262676 -5156 262678
rect 589080 262676 589680 262678
rect -5756 262074 -5156 262076
rect 589080 262074 589680 262076
rect 0 259396 584000 261756
rect -3876 259076 -3276 259078
rect 587200 259076 587800 259078
rect -3876 258474 -3276 258476
rect 587200 258474 587800 258476
rect 0 255748 584000 258156
rect -1996 255428 -1396 255430
rect 585320 255428 585920 255430
rect -1996 254826 -1396 254828
rect 585320 254826 585920 254828
rect 0 248596 584000 254508
rect -8576 248276 -7976 248278
rect 591900 248276 592500 248278
rect -8576 247674 -7976 247676
rect 591900 247674 592500 247676
rect 0 244996 584000 247356
rect -6696 244676 -6096 244678
rect 590020 244676 590620 244678
rect -6696 244074 -6096 244076
rect 590020 244074 590620 244076
rect 0 241396 584000 243756
rect -4816 241076 -4216 241078
rect 588140 241076 588740 241078
rect -4816 240474 -4216 240476
rect 588140 240474 588740 240476
rect 0 237748 584000 240156
rect -2936 237428 -2336 237430
rect 586260 237428 586860 237430
rect -2936 236826 -2336 236828
rect 586260 236826 586860 236828
rect 0 230596 584000 236508
rect -7636 230276 -7036 230278
rect 590960 230276 591560 230278
rect -7636 229674 -7036 229676
rect 590960 229674 591560 229676
rect 0 226996 584000 229356
rect -5756 226676 -5156 226678
rect 589080 226676 589680 226678
rect -5756 226074 -5156 226076
rect 589080 226074 589680 226076
rect 0 223396 584000 225756
rect -3876 223076 -3276 223078
rect 587200 223076 587800 223078
rect -3876 222474 -3276 222476
rect 587200 222474 587800 222476
rect 0 219748 584000 222156
rect -1996 219428 -1396 219430
rect 585320 219428 585920 219430
rect -1996 218826 -1396 218828
rect 585320 218826 585920 218828
rect 0 212596 584000 218508
rect -8576 212276 -7976 212278
rect 591900 212276 592500 212278
rect -8576 211674 -7976 211676
rect 591900 211674 592500 211676
rect 0 208996 584000 211356
rect -6696 208676 -6096 208678
rect 590020 208676 590620 208678
rect -6696 208074 -6096 208076
rect 590020 208074 590620 208076
rect 0 205396 584000 207756
rect -4816 205076 -4216 205078
rect 588140 205076 588740 205078
rect -4816 204474 -4216 204476
rect 588140 204474 588740 204476
rect 0 201748 584000 204156
rect -2936 201428 -2336 201430
rect 586260 201428 586860 201430
rect -2936 200826 -2336 200828
rect 586260 200826 586860 200828
rect 0 194596 584000 200508
rect -7636 194276 -7036 194278
rect 590960 194276 591560 194278
rect -7636 193674 -7036 193676
rect 590960 193674 591560 193676
rect 0 190996 584000 193356
rect -5756 190676 -5156 190678
rect 589080 190676 589680 190678
rect -5756 190074 -5156 190076
rect 589080 190074 589680 190076
rect 0 187396 584000 189756
rect -3876 187076 -3276 187078
rect 587200 187076 587800 187078
rect -3876 186474 -3276 186476
rect 587200 186474 587800 186476
rect 0 183748 584000 186156
rect -1996 183428 -1396 183430
rect 585320 183428 585920 183430
rect -1996 182826 -1396 182828
rect 585320 182826 585920 182828
rect 0 176596 584000 182508
rect -8576 176276 -7976 176278
rect 591900 176276 592500 176278
rect -8576 175674 -7976 175676
rect 591900 175674 592500 175676
rect 0 172996 584000 175356
rect -6696 172676 -6096 172678
rect 590020 172676 590620 172678
rect -6696 172074 -6096 172076
rect 590020 172074 590620 172076
rect 0 169396 584000 171756
rect -4816 169076 -4216 169078
rect 588140 169076 588740 169078
rect -4816 168474 -4216 168476
rect 588140 168474 588740 168476
rect 0 165748 584000 168156
rect -2936 165428 -2336 165430
rect 586260 165428 586860 165430
rect -2936 164826 -2336 164828
rect 586260 164826 586860 164828
rect 0 158596 584000 164508
rect -7636 158276 -7036 158278
rect 590960 158276 591560 158278
rect -7636 157674 -7036 157676
rect 590960 157674 591560 157676
rect 0 154996 584000 157356
rect -5756 154676 -5156 154678
rect 589080 154676 589680 154678
rect -5756 154074 -5156 154076
rect 589080 154074 589680 154076
rect 0 151396 584000 153756
rect -3876 151076 -3276 151078
rect 587200 151076 587800 151078
rect -3876 150474 -3276 150476
rect 587200 150474 587800 150476
rect 0 147748 584000 150156
rect -1996 147428 -1396 147430
rect 585320 147428 585920 147430
rect -1996 146826 -1396 146828
rect 585320 146826 585920 146828
rect 0 140596 584000 146508
rect -8576 140276 -7976 140278
rect 591900 140276 592500 140278
rect -8576 139674 -7976 139676
rect 591900 139674 592500 139676
rect 0 136996 584000 139356
rect -6696 136676 -6096 136678
rect 590020 136676 590620 136678
rect -6696 136074 -6096 136076
rect 590020 136074 590620 136076
rect 0 133396 584000 135756
rect -4816 133076 -4216 133078
rect 588140 133076 588740 133078
rect -4816 132474 -4216 132476
rect 588140 132474 588740 132476
rect 0 129748 584000 132156
rect -2936 129428 -2336 129430
rect 586260 129428 586860 129430
rect -2936 128826 -2336 128828
rect 586260 128826 586860 128828
rect 0 122596 584000 128508
rect -7636 122276 -7036 122278
rect 590960 122276 591560 122278
rect -7636 121674 -7036 121676
rect 590960 121674 591560 121676
rect 0 118996 584000 121356
rect -5756 118676 -5156 118678
rect 589080 118676 589680 118678
rect -5756 118074 -5156 118076
rect 589080 118074 589680 118076
rect 0 115396 584000 117756
rect -3876 115076 -3276 115078
rect 587200 115076 587800 115078
rect -3876 114474 -3276 114476
rect 587200 114474 587800 114476
rect 0 111748 584000 114156
rect -1996 111428 -1396 111430
rect 585320 111428 585920 111430
rect -1996 110826 -1396 110828
rect 585320 110826 585920 110828
rect 0 104596 584000 110508
rect -8576 104276 -7976 104278
rect 591900 104276 592500 104278
rect -8576 103674 -7976 103676
rect 591900 103674 592500 103676
rect 0 100996 584000 103356
rect -6696 100676 -6096 100678
rect 590020 100676 590620 100678
rect -6696 100074 -6096 100076
rect 590020 100074 590620 100076
rect 0 97396 584000 99756
rect -4816 97076 -4216 97078
rect 588140 97076 588740 97078
rect -4816 96474 -4216 96476
rect 588140 96474 588740 96476
rect 0 93748 584000 96156
rect -2936 93428 -2336 93430
rect 586260 93428 586860 93430
rect -2936 92826 -2336 92828
rect 586260 92826 586860 92828
rect 0 86596 584000 92508
rect -7636 86276 -7036 86278
rect 590960 86276 591560 86278
rect -7636 85674 -7036 85676
rect 590960 85674 591560 85676
rect 0 82996 584000 85356
rect -5756 82676 -5156 82678
rect 589080 82676 589680 82678
rect -5756 82074 -5156 82076
rect 589080 82074 589680 82076
rect 0 79396 584000 81756
rect -3876 79076 -3276 79078
rect 587200 79076 587800 79078
rect -3876 78474 -3276 78476
rect 587200 78474 587800 78476
rect 0 75748 584000 78156
rect -1996 75428 -1396 75430
rect 585320 75428 585920 75430
rect -1996 74826 -1396 74828
rect 585320 74826 585920 74828
rect 0 68596 584000 74508
rect -8576 68276 -7976 68278
rect 591900 68276 592500 68278
rect -8576 67674 -7976 67676
rect 591900 67674 592500 67676
rect 0 64996 584000 67356
rect -6696 64676 -6096 64678
rect 590020 64676 590620 64678
rect -6696 64074 -6096 64076
rect 590020 64074 590620 64076
rect 0 61396 584000 63756
rect -4816 61076 -4216 61078
rect 588140 61076 588740 61078
rect -4816 60474 -4216 60476
rect 588140 60474 588740 60476
rect 0 57748 584000 60156
rect -2936 57428 -2336 57430
rect 586260 57428 586860 57430
rect -2936 56826 -2336 56828
rect 586260 56826 586860 56828
rect 0 50596 584000 56508
rect -7636 50276 -7036 50278
rect 590960 50276 591560 50278
rect -7636 49674 -7036 49676
rect 590960 49674 591560 49676
rect 0 46996 584000 49356
rect -5756 46676 -5156 46678
rect 589080 46676 589680 46678
rect -5756 46074 -5156 46076
rect 589080 46074 589680 46076
rect 0 43396 584000 45756
rect -3876 43076 -3276 43078
rect 587200 43076 587800 43078
rect -3876 42474 -3276 42476
rect 587200 42474 587800 42476
rect 0 39748 584000 42156
rect -1996 39428 -1396 39430
rect 585320 39428 585920 39430
rect -1996 38826 -1396 38828
rect 585320 38826 585920 38828
rect 0 32596 584000 38508
rect -8576 32276 -7976 32278
rect 591900 32276 592500 32278
rect -8576 31674 -7976 31676
rect 591900 31674 592500 31676
rect 0 28996 584000 31356
rect -6696 28676 -6096 28678
rect 590020 28676 590620 28678
rect -6696 28074 -6096 28076
rect 590020 28074 590620 28076
rect 0 25396 584000 27756
rect -4816 25076 -4216 25078
rect 588140 25076 588740 25078
rect -4816 24474 -4216 24476
rect 588140 24474 588740 24476
rect 0 21748 584000 24156
rect -2936 21428 -2336 21430
rect 586260 21428 586860 21430
rect -2936 20826 -2336 20828
rect 586260 20826 586860 20828
rect 0 14596 584000 20508
rect -7636 14276 -7036 14278
rect 590960 14276 591560 14278
rect -7636 13674 -7036 13676
rect 590960 13674 591560 13676
rect 0 10996 584000 13356
rect -5756 10676 -5156 10678
rect 589080 10676 589680 10678
rect -5756 10074 -5156 10076
rect 589080 10074 589680 10076
rect 0 7396 584000 9756
rect -3876 7076 -3276 7078
rect 587200 7076 587800 7078
rect -3876 6474 -3276 6476
rect 587200 6474 587800 6476
rect 0 3748 584000 6156
rect -1996 3428 -1396 3430
rect 585320 3428 585920 3430
rect -1996 2826 -1396 2828
rect 585320 2826 585920 2828
rect 0 0 584000 2508
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
<< labels >>
rlabel metal3 s 583520 5660 584960 5900 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 467244 584960 467484 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 513348 584960 513588 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 559452 584960 559692 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 605692 584960 605932 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 583520 651796 584960 652036 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 576830 703520 576942 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 519790 703520 519902 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 462842 703520 462954 704960 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 405894 703520 406006 704960 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 348854 703520 348966 704960 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 51764 584960 52004 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 291906 703520 292018 704960 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 234958 703520 235070 704960 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 177918 703520 178030 704960 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 120970 703520 121082 704960 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 697628 480 697868 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 648124 480 648364 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 598756 480 598996 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 549388 480 549628 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 500020 480 500260 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s -960 450652 480 450892 4 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 97868 584960 98108 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s -960 401148 480 401388 4 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 698036 584960 698276 6 analog_io[31]
port 25 nsew signal bidirectional
rlabel metal2 s 64022 703520 64134 704960 6 analog_io[32]
port 26 nsew signal bidirectional
rlabel metal2 s 49762 703520 49874 704960 6 analog_io[33]
port 27 nsew signal bidirectional
rlabel metal3 s -960 92428 480 92668 4 analog_io[34]
port 28 nsew signal bidirectional
rlabel metal2 s 577474 -960 577586 480 8 analog_io[35]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 144108 584960 144348 6 analog_io[3]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 190212 584960 190452 6 analog_io[4]
port 31 nsew signal bidirectional
rlabel metal3 s 583520 236452 584960 236692 6 analog_io[5]
port 32 nsew signal bidirectional
rlabel metal3 s 583520 282556 584960 282796 6 analog_io[6]
port 33 nsew signal bidirectional
rlabel metal3 s 583520 328660 584960 328900 6 analog_io[7]
port 34 nsew signal bidirectional
rlabel metal3 s 583520 374900 584960 375140 6 analog_io[8]
port 35 nsew signal bidirectional
rlabel metal3 s 583520 421004 584960 421244 6 analog_io[9]
port 36 nsew signal bidirectional
rlabel metal3 s 583520 17084 584960 17324 6 io_in[0]
port 37 nsew signal input
rlabel metal3 s 583520 478668 584960 478908 6 io_in[10]
port 38 nsew signal input
rlabel metal3 s 583520 524908 584960 525148 6 io_in[11]
port 39 nsew signal input
rlabel metal3 s 583520 571012 584960 571252 6 io_in[12]
port 40 nsew signal input
rlabel metal3 s 583520 617252 584960 617492 6 io_in[13]
port 41 nsew signal input
rlabel metal3 s 583520 663356 584960 663596 6 io_in[14]
port 42 nsew signal input
rlabel metal2 s 562570 703520 562682 704960 6 io_in[15]
port 43 nsew signal input
rlabel metal2 s 505622 703520 505734 704960 6 io_in[16]
port 44 nsew signal input
rlabel metal2 s 448582 703520 448694 704960 6 io_in[17]
port 45 nsew signal input
rlabel metal2 s 391634 703520 391746 704960 6 io_in[18]
port 46 nsew signal input
rlabel metal2 s 334686 703520 334798 704960 6 io_in[19]
port 47 nsew signal input
rlabel metal3 s 583520 63324 584960 63564 6 io_in[1]
port 48 nsew signal input
rlabel metal2 s 277646 703520 277758 704960 6 io_in[20]
port 49 nsew signal input
rlabel metal2 s 220698 703520 220810 704960 6 io_in[21]
port 50 nsew signal input
rlabel metal2 s 163750 703520 163862 704960 6 io_in[22]
port 51 nsew signal input
rlabel metal2 s 106710 703520 106822 704960 6 io_in[23]
port 52 nsew signal input
rlabel metal3 s -960 685252 480 685492 4 io_in[24]
port 53 nsew signal input
rlabel metal3 s -960 635884 480 636124 4 io_in[25]
port 54 nsew signal input
rlabel metal3 s -960 586380 480 586620 4 io_in[26]
port 55 nsew signal input
rlabel metal3 s -960 537012 480 537252 4 io_in[27]
port 56 nsew signal input
rlabel metal3 s -960 487644 480 487884 4 io_in[28]
port 57 nsew signal input
rlabel metal3 s -960 438276 480 438516 4 io_in[29]
port 58 nsew signal input
rlabel metal3 s 583520 109428 584960 109668 6 io_in[2]
port 59 nsew signal input
rlabel metal3 s -960 388908 480 389148 4 io_in[30]
port 60 nsew signal input
rlabel metal3 s -960 351780 480 352020 4 io_in[31]
port 61 nsew signal input
rlabel metal3 s -960 314788 480 315028 4 io_in[32]
port 62 nsew signal input
rlabel metal3 s -960 277660 480 277900 4 io_in[33]
port 63 nsew signal input
rlabel metal3 s -960 240668 480 240908 4 io_in[34]
port 64 nsew signal input
rlabel metal3 s -960 203540 480 203780 4 io_in[35]
port 65 nsew signal input
rlabel metal3 s -960 166548 480 166788 4 io_in[36]
port 66 nsew signal input
rlabel metal3 s -960 129556 480 129796 4 io_in[37]
port 67 nsew signal input
rlabel metal2 s 578670 -960 578782 480 8 io_in[38]
port 68 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 io_in[39]
port 69 nsew signal input
rlabel metal3 s 583520 155668 584960 155908 6 io_in[3]
port 70 nsew signal input
rlabel metal2 s 21242 703520 21354 704960 6 io_in[40]
port 71 nsew signal input
rlabel metal3 s -960 30684 480 30924 4 io_in[41]
port 72 nsew signal input
rlabel metal2 s 7074 703520 7186 704960 6 io_in[42]
port 73 nsew signal input
rlabel metal3 s 583520 201772 584960 202012 6 io_in[4]
port 74 nsew signal input
rlabel metal3 s 583520 247876 584960 248116 6 io_in[5]
port 75 nsew signal input
rlabel metal3 s 583520 294116 584960 294356 6 io_in[6]
port 76 nsew signal input
rlabel metal3 s 583520 340220 584960 340460 6 io_in[7]
port 77 nsew signal input
rlabel metal3 s 583520 386460 584960 386700 6 io_in[8]
port 78 nsew signal input
rlabel metal3 s 583520 432564 584960 432804 6 io_in[9]
port 79 nsew signal input
rlabel metal3 s 583520 40204 584960 40444 6 io_oeb[0]
port 80 nsew signal output
rlabel metal3 s 583520 501788 584960 502028 6 io_oeb[10]
port 81 nsew signal output
rlabel metal3 s 583520 548028 584960 548268 6 io_oeb[11]
port 82 nsew signal output
rlabel metal3 s 583520 594132 584960 594372 6 io_oeb[12]
port 83 nsew signal output
rlabel metal3 s 583520 640236 584960 640476 6 io_oeb[13]
port 84 nsew signal output
rlabel metal3 s 583520 686476 584960 686716 6 io_oeb[14]
port 85 nsew signal output
rlabel metal2 s 534050 703520 534162 704960 6 io_oeb[15]
port 86 nsew signal output
rlabel metal2 s 477102 703520 477214 704960 6 io_oeb[16]
port 87 nsew signal output
rlabel metal2 s 420154 703520 420266 704960 6 io_oeb[17]
port 88 nsew signal output
rlabel metal2 s 363114 703520 363226 704960 6 io_oeb[18]
port 89 nsew signal output
rlabel metal2 s 306166 703520 306278 704960 6 io_oeb[19]
port 90 nsew signal output
rlabel metal3 s 583520 86308 584960 86548 6 io_oeb[1]
port 91 nsew signal output
rlabel metal2 s 249218 703520 249330 704960 6 io_oeb[20]
port 92 nsew signal output
rlabel metal2 s 192178 703520 192290 704960 6 io_oeb[21]
port 93 nsew signal output
rlabel metal2 s 135230 703520 135342 704960 6 io_oeb[22]
port 94 nsew signal output
rlabel metal2 s 78282 703520 78394 704960 6 io_oeb[23]
port 95 nsew signal output
rlabel metal3 s -960 660500 480 660740 4 io_oeb[24]
port 96 nsew signal output
rlabel metal3 s -960 611132 480 611372 4 io_oeb[25]
port 97 nsew signal output
rlabel metal3 s -960 561764 480 562004 4 io_oeb[26]
port 98 nsew signal output
rlabel metal3 s -960 512396 480 512636 4 io_oeb[27]
port 99 nsew signal output
rlabel metal3 s -960 462892 480 463132 4 io_oeb[28]
port 100 nsew signal output
rlabel metal3 s -960 413524 480 413764 4 io_oeb[29]
port 101 nsew signal output
rlabel metal3 s 583520 132548 584960 132788 6 io_oeb[2]
port 102 nsew signal output
rlabel metal3 s -960 364156 480 364396 4 io_oeb[30]
port 103 nsew signal output
rlabel metal3 s -960 327028 480 327268 4 io_oeb[31]
port 104 nsew signal output
rlabel metal3 s -960 290036 480 290276 4 io_oeb[32]
port 105 nsew signal output
rlabel metal3 s -960 253044 480 253284 4 io_oeb[33]
port 106 nsew signal output
rlabel metal3 s -960 215916 480 216156 4 io_oeb[34]
port 107 nsew signal output
rlabel metal3 s -960 178924 480 179164 4 io_oeb[35]
port 108 nsew signal output
rlabel metal3 s -960 141796 480 142036 4 io_oeb[36]
port 109 nsew signal output
rlabel metal3 s -960 104804 480 105044 4 io_oeb[37]
port 110 nsew signal output
rlabel metal3 s -960 80052 480 80292 4 io_oeb[38]
port 111 nsew signal output
rlabel metal3 s -960 55436 480 55676 4 io_oeb[39]
port 112 nsew signal output
rlabel metal3 s 583520 178652 584960 178892 6 io_oeb[3]
port 113 nsew signal output
rlabel metal3 s -960 43060 480 43300 4 io_oeb[40]
port 114 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 io_oeb[41]
port 115 nsew signal output
rlabel metal3 s -960 18308 480 18548 4 io_oeb[42]
port 116 nsew signal output
rlabel metal3 s 583520 224892 584960 225132 6 io_oeb[4]
port 117 nsew signal output
rlabel metal3 s 583520 270996 584960 271236 6 io_oeb[5]
port 118 nsew signal output
rlabel metal3 s 583520 317236 584960 317476 6 io_oeb[6]
port 119 nsew signal output
rlabel metal3 s 583520 363340 584960 363580 6 io_oeb[7]
port 120 nsew signal output
rlabel metal3 s 583520 409444 584960 409684 6 io_oeb[8]
port 121 nsew signal output
rlabel metal3 s 583520 455684 584960 455924 6 io_oeb[9]
port 122 nsew signal output
rlabel metal3 s 583520 28644 584960 28884 6 io_out[0]
port 123 nsew signal output
rlabel metal3 s 583520 490228 584960 490468 6 io_out[10]
port 124 nsew signal output
rlabel metal3 s 583520 536468 584960 536708 6 io_out[11]
port 125 nsew signal output
rlabel metal3 s 583520 582572 584960 582812 6 io_out[12]
port 126 nsew signal output
rlabel metal3 s 583520 628812 584960 629052 6 io_out[13]
port 127 nsew signal output
rlabel metal3 s 583520 674916 584960 675156 6 io_out[14]
port 128 nsew signal output
rlabel metal2 s 548310 703520 548422 704960 6 io_out[15]
port 129 nsew signal output
rlabel metal2 s 491362 703520 491474 704960 6 io_out[16]
port 130 nsew signal output
rlabel metal2 s 434322 703520 434434 704960 6 io_out[17]
port 131 nsew signal output
rlabel metal2 s 377374 703520 377486 704960 6 io_out[18]
port 132 nsew signal output
rlabel metal2 s 320426 703520 320538 704960 6 io_out[19]
port 133 nsew signal output
rlabel metal3 s 583520 74884 584960 75124 6 io_out[1]
port 134 nsew signal output
rlabel metal2 s 263386 703520 263498 704960 6 io_out[20]
port 135 nsew signal output
rlabel metal2 s 206438 703520 206550 704960 6 io_out[21]
port 136 nsew signal output
rlabel metal2 s 149490 703520 149602 704960 6 io_out[22]
port 137 nsew signal output
rlabel metal2 s 92450 703520 92562 704960 6 io_out[23]
port 138 nsew signal output
rlabel metal3 s -960 672876 480 673116 4 io_out[24]
port 139 nsew signal output
rlabel metal3 s -960 623508 480 623748 4 io_out[25]
port 140 nsew signal output
rlabel metal3 s -960 574140 480 574380 4 io_out[26]
port 141 nsew signal output
rlabel metal3 s -960 524636 480 524876 4 io_out[27]
port 142 nsew signal output
rlabel metal3 s -960 475268 480 475508 4 io_out[28]
port 143 nsew signal output
rlabel metal3 s -960 425900 480 426140 4 io_out[29]
port 144 nsew signal output
rlabel metal3 s 583520 120988 584960 121228 6 io_out[2]
port 145 nsew signal output
rlabel metal3 s -960 376532 480 376772 4 io_out[30]
port 146 nsew signal output
rlabel metal3 s -960 339404 480 339644 4 io_out[31]
port 147 nsew signal output
rlabel metal3 s -960 302412 480 302652 4 io_out[32]
port 148 nsew signal output
rlabel metal3 s -960 265284 480 265524 4 io_out[33]
port 149 nsew signal output
rlabel metal3 s -960 228292 480 228532 4 io_out[34]
port 150 nsew signal output
rlabel metal3 s -960 191300 480 191540 4 io_out[35]
port 151 nsew signal output
rlabel metal3 s -960 154172 480 154412 4 io_out[36]
port 152 nsew signal output
rlabel metal3 s -960 117180 480 117420 4 io_out[37]
port 153 nsew signal output
rlabel metal3 s -960 67812 480 68052 4 io_out[38]
port 154 nsew signal output
rlabel metal2 s 35502 703520 35614 704960 6 io_out[39]
port 155 nsew signal output
rlabel metal3 s 583520 167092 584960 167332 6 io_out[3]
port 156 nsew signal output
rlabel metal2 s 580970 -960 581082 480 8 io_out[40]
port 157 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 io_out[41]
port 158 nsew signal output
rlabel metal3 s -960 6068 480 6308 4 io_out[42]
port 159 nsew signal output
rlabel metal3 s 583520 213332 584960 213572 6 io_out[4]
port 160 nsew signal output
rlabel metal3 s 583520 259436 584960 259676 6 io_out[5]
port 161 nsew signal output
rlabel metal3 s 583520 305676 584960 305916 6 io_out[6]
port 162 nsew signal output
rlabel metal3 s 583520 351780 584960 352020 6 io_out[7]
port 163 nsew signal output
rlabel metal3 s 583520 397884 584960 398124 6 io_out[8]
port 164 nsew signal output
rlabel metal3 s 583520 444124 584960 444364 6 io_out[9]
port 165 nsew signal output
rlabel metal2 s 125018 -960 125130 480 8 la_data_in[0]
port 166 nsew signal input
rlabel metal2 s 477562 -960 477674 480 8 la_data_in[100]
port 167 nsew signal input
rlabel metal2 s 481150 -960 481262 480 8 la_data_in[101]
port 168 nsew signal input
rlabel metal2 s 484646 -960 484758 480 8 la_data_in[102]
port 169 nsew signal input
rlabel metal2 s 488142 -960 488254 480 8 la_data_in[103]
port 170 nsew signal input
rlabel metal2 s 491638 -960 491750 480 8 la_data_in[104]
port 171 nsew signal input
rlabel metal2 s 495226 -960 495338 480 8 la_data_in[105]
port 172 nsew signal input
rlabel metal2 s 498722 -960 498834 480 8 la_data_in[106]
port 173 nsew signal input
rlabel metal2 s 502218 -960 502330 480 8 la_data_in[107]
port 174 nsew signal input
rlabel metal2 s 505806 -960 505918 480 8 la_data_in[108]
port 175 nsew signal input
rlabel metal2 s 509302 -960 509414 480 8 la_data_in[109]
port 176 nsew signal input
rlabel metal2 s 160346 -960 160458 480 8 la_data_in[10]
port 177 nsew signal input
rlabel metal2 s 512798 -960 512910 480 8 la_data_in[110]
port 178 nsew signal input
rlabel metal2 s 516386 -960 516498 480 8 la_data_in[111]
port 179 nsew signal input
rlabel metal2 s 519882 -960 519994 480 8 la_data_in[112]
port 180 nsew signal input
rlabel metal2 s 523378 -960 523490 480 8 la_data_in[113]
port 181 nsew signal input
rlabel metal2 s 526966 -960 527078 480 8 la_data_in[114]
port 182 nsew signal input
rlabel metal2 s 530462 -960 530574 480 8 la_data_in[115]
port 183 nsew signal input
rlabel metal2 s 533958 -960 534070 480 8 la_data_in[116]
port 184 nsew signal input
rlabel metal2 s 537546 -960 537658 480 8 la_data_in[117]
port 185 nsew signal input
rlabel metal2 s 541042 -960 541154 480 8 la_data_in[118]
port 186 nsew signal input
rlabel metal2 s 544538 -960 544650 480 8 la_data_in[119]
port 187 nsew signal input
rlabel metal2 s 163842 -960 163954 480 8 la_data_in[11]
port 188 nsew signal input
rlabel metal2 s 548126 -960 548238 480 8 la_data_in[120]
port 189 nsew signal input
rlabel metal2 s 551622 -960 551734 480 8 la_data_in[121]
port 190 nsew signal input
rlabel metal2 s 555118 -960 555230 480 8 la_data_in[122]
port 191 nsew signal input
rlabel metal2 s 558706 -960 558818 480 8 la_data_in[123]
port 192 nsew signal input
rlabel metal2 s 562202 -960 562314 480 8 la_data_in[124]
port 193 nsew signal input
rlabel metal2 s 565698 -960 565810 480 8 la_data_in[125]
port 194 nsew signal input
rlabel metal2 s 569194 -960 569306 480 8 la_data_in[126]
port 195 nsew signal input
rlabel metal2 s 572782 -960 572894 480 8 la_data_in[127]
port 196 nsew signal input
rlabel metal2 s 167338 -960 167450 480 8 la_data_in[12]
port 197 nsew signal input
rlabel metal2 s 170926 -960 171038 480 8 la_data_in[13]
port 198 nsew signal input
rlabel metal2 s 174422 -960 174534 480 8 la_data_in[14]
port 199 nsew signal input
rlabel metal2 s 177918 -960 178030 480 8 la_data_in[15]
port 200 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_data_in[16]
port 201 nsew signal input
rlabel metal2 s 185002 -960 185114 480 8 la_data_in[17]
port 202 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_data_in[18]
port 203 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_data_in[19]
port 204 nsew signal input
rlabel metal2 s 128606 -960 128718 480 8 la_data_in[1]
port 205 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_data_in[20]
port 206 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_data_in[21]
port 207 nsew signal input
rlabel metal2 s 202574 -960 202686 480 8 la_data_in[22]
port 208 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_data_in[23]
port 209 nsew signal input
rlabel metal2 s 209658 -960 209770 480 8 la_data_in[24]
port 210 nsew signal input
rlabel metal2 s 213154 -960 213266 480 8 la_data_in[25]
port 211 nsew signal input
rlabel metal2 s 216742 -960 216854 480 8 la_data_in[26]
port 212 nsew signal input
rlabel metal2 s 220238 -960 220350 480 8 la_data_in[27]
port 213 nsew signal input
rlabel metal2 s 223734 -960 223846 480 8 la_data_in[28]
port 214 nsew signal input
rlabel metal2 s 227322 -960 227434 480 8 la_data_in[29]
port 215 nsew signal input
rlabel metal2 s 132102 -960 132214 480 8 la_data_in[2]
port 216 nsew signal input
rlabel metal2 s 230818 -960 230930 480 8 la_data_in[30]
port 217 nsew signal input
rlabel metal2 s 234314 -960 234426 480 8 la_data_in[31]
port 218 nsew signal input
rlabel metal2 s 237902 -960 238014 480 8 la_data_in[32]
port 219 nsew signal input
rlabel metal2 s 241398 -960 241510 480 8 la_data_in[33]
port 220 nsew signal input
rlabel metal2 s 244894 -960 245006 480 8 la_data_in[34]
port 221 nsew signal input
rlabel metal2 s 248482 -960 248594 480 8 la_data_in[35]
port 222 nsew signal input
rlabel metal2 s 251978 -960 252090 480 8 la_data_in[36]
port 223 nsew signal input
rlabel metal2 s 255474 -960 255586 480 8 la_data_in[37]
port 224 nsew signal input
rlabel metal2 s 258970 -960 259082 480 8 la_data_in[38]
port 225 nsew signal input
rlabel metal2 s 262558 -960 262670 480 8 la_data_in[39]
port 226 nsew signal input
rlabel metal2 s 135598 -960 135710 480 8 la_data_in[3]
port 227 nsew signal input
rlabel metal2 s 266054 -960 266166 480 8 la_data_in[40]
port 228 nsew signal input
rlabel metal2 s 269550 -960 269662 480 8 la_data_in[41]
port 229 nsew signal input
rlabel metal2 s 273138 -960 273250 480 8 la_data_in[42]
port 230 nsew signal input
rlabel metal2 s 276634 -960 276746 480 8 la_data_in[43]
port 231 nsew signal input
rlabel metal2 s 280130 -960 280242 480 8 la_data_in[44]
port 232 nsew signal input
rlabel metal2 s 283718 -960 283830 480 8 la_data_in[45]
port 233 nsew signal input
rlabel metal2 s 287214 -960 287326 480 8 la_data_in[46]
port 234 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[47]
port 235 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[48]
port 236 nsew signal input
rlabel metal2 s 297794 -960 297906 480 8 la_data_in[49]
port 237 nsew signal input
rlabel metal2 s 139186 -960 139298 480 8 la_data_in[4]
port 238 nsew signal input
rlabel metal2 s 301290 -960 301402 480 8 la_data_in[50]
port 239 nsew signal input
rlabel metal2 s 304878 -960 304990 480 8 la_data_in[51]
port 240 nsew signal input
rlabel metal2 s 308374 -960 308486 480 8 la_data_in[52]
port 241 nsew signal input
rlabel metal2 s 311870 -960 311982 480 8 la_data_in[53]
port 242 nsew signal input
rlabel metal2 s 315458 -960 315570 480 8 la_data_in[54]
port 243 nsew signal input
rlabel metal2 s 318954 -960 319066 480 8 la_data_in[55]
port 244 nsew signal input
rlabel metal2 s 322450 -960 322562 480 8 la_data_in[56]
port 245 nsew signal input
rlabel metal2 s 326038 -960 326150 480 8 la_data_in[57]
port 246 nsew signal input
rlabel metal2 s 329534 -960 329646 480 8 la_data_in[58]
port 247 nsew signal input
rlabel metal2 s 333030 -960 333142 480 8 la_data_in[59]
port 248 nsew signal input
rlabel metal2 s 142682 -960 142794 480 8 la_data_in[5]
port 249 nsew signal input
rlabel metal2 s 336526 -960 336638 480 8 la_data_in[60]
port 250 nsew signal input
rlabel metal2 s 340114 -960 340226 480 8 la_data_in[61]
port 251 nsew signal input
rlabel metal2 s 343610 -960 343722 480 8 la_data_in[62]
port 252 nsew signal input
rlabel metal2 s 347106 -960 347218 480 8 la_data_in[63]
port 253 nsew signal input
rlabel metal2 s 350694 -960 350806 480 8 la_data_in[64]
port 254 nsew signal input
rlabel metal2 s 354190 -960 354302 480 8 la_data_in[65]
port 255 nsew signal input
rlabel metal2 s 357686 -960 357798 480 8 la_data_in[66]
port 256 nsew signal input
rlabel metal2 s 361274 -960 361386 480 8 la_data_in[67]
port 257 nsew signal input
rlabel metal2 s 364770 -960 364882 480 8 la_data_in[68]
port 258 nsew signal input
rlabel metal2 s 368266 -960 368378 480 8 la_data_in[69]
port 259 nsew signal input
rlabel metal2 s 146178 -960 146290 480 8 la_data_in[6]
port 260 nsew signal input
rlabel metal2 s 371854 -960 371966 480 8 la_data_in[70]
port 261 nsew signal input
rlabel metal2 s 375350 -960 375462 480 8 la_data_in[71]
port 262 nsew signal input
rlabel metal2 s 378846 -960 378958 480 8 la_data_in[72]
port 263 nsew signal input
rlabel metal2 s 382434 -960 382546 480 8 la_data_in[73]
port 264 nsew signal input
rlabel metal2 s 385930 -960 386042 480 8 la_data_in[74]
port 265 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_data_in[75]
port 266 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_data_in[76]
port 267 nsew signal input
rlabel metal2 s 396510 -960 396622 480 8 la_data_in[77]
port 268 nsew signal input
rlabel metal2 s 400006 -960 400118 480 8 la_data_in[78]
port 269 nsew signal input
rlabel metal2 s 403594 -960 403706 480 8 la_data_in[79]
port 270 nsew signal input
rlabel metal2 s 149766 -960 149878 480 8 la_data_in[7]
port 271 nsew signal input
rlabel metal2 s 407090 -960 407202 480 8 la_data_in[80]
port 272 nsew signal input
rlabel metal2 s 410586 -960 410698 480 8 la_data_in[81]
port 273 nsew signal input
rlabel metal2 s 414082 -960 414194 480 8 la_data_in[82]
port 274 nsew signal input
rlabel metal2 s 417670 -960 417782 480 8 la_data_in[83]
port 275 nsew signal input
rlabel metal2 s 421166 -960 421278 480 8 la_data_in[84]
port 276 nsew signal input
rlabel metal2 s 424662 -960 424774 480 8 la_data_in[85]
port 277 nsew signal input
rlabel metal2 s 428250 -960 428362 480 8 la_data_in[86]
port 278 nsew signal input
rlabel metal2 s 431746 -960 431858 480 8 la_data_in[87]
port 279 nsew signal input
rlabel metal2 s 435242 -960 435354 480 8 la_data_in[88]
port 280 nsew signal input
rlabel metal2 s 438830 -960 438942 480 8 la_data_in[89]
port 281 nsew signal input
rlabel metal2 s 153262 -960 153374 480 8 la_data_in[8]
port 282 nsew signal input
rlabel metal2 s 442326 -960 442438 480 8 la_data_in[90]
port 283 nsew signal input
rlabel metal2 s 445822 -960 445934 480 8 la_data_in[91]
port 284 nsew signal input
rlabel metal2 s 449410 -960 449522 480 8 la_data_in[92]
port 285 nsew signal input
rlabel metal2 s 452906 -960 453018 480 8 la_data_in[93]
port 286 nsew signal input
rlabel metal2 s 456402 -960 456514 480 8 la_data_in[94]
port 287 nsew signal input
rlabel metal2 s 459990 -960 460102 480 8 la_data_in[95]
port 288 nsew signal input
rlabel metal2 s 463486 -960 463598 480 8 la_data_in[96]
port 289 nsew signal input
rlabel metal2 s 466982 -960 467094 480 8 la_data_in[97]
port 290 nsew signal input
rlabel metal2 s 470570 -960 470682 480 8 la_data_in[98]
port 291 nsew signal input
rlabel metal2 s 474066 -960 474178 480 8 la_data_in[99]
port 292 nsew signal input
rlabel metal2 s 156758 -960 156870 480 8 la_data_in[9]
port 293 nsew signal input
rlabel metal2 s 126214 -960 126326 480 8 la_data_out[0]
port 294 nsew signal output
rlabel metal2 s 478758 -960 478870 480 8 la_data_out[100]
port 295 nsew signal output
rlabel metal2 s 482254 -960 482366 480 8 la_data_out[101]
port 296 nsew signal output
rlabel metal2 s 485842 -960 485954 480 8 la_data_out[102]
port 297 nsew signal output
rlabel metal2 s 489338 -960 489450 480 8 la_data_out[103]
port 298 nsew signal output
rlabel metal2 s 492834 -960 492946 480 8 la_data_out[104]
port 299 nsew signal output
rlabel metal2 s 496422 -960 496534 480 8 la_data_out[105]
port 300 nsew signal output
rlabel metal2 s 499918 -960 500030 480 8 la_data_out[106]
port 301 nsew signal output
rlabel metal2 s 503414 -960 503526 480 8 la_data_out[107]
port 302 nsew signal output
rlabel metal2 s 507002 -960 507114 480 8 la_data_out[108]
port 303 nsew signal output
rlabel metal2 s 510498 -960 510610 480 8 la_data_out[109]
port 304 nsew signal output
rlabel metal2 s 161450 -960 161562 480 8 la_data_out[10]
port 305 nsew signal output
rlabel metal2 s 513994 -960 514106 480 8 la_data_out[110]
port 306 nsew signal output
rlabel metal2 s 517490 -960 517602 480 8 la_data_out[111]
port 307 nsew signal output
rlabel metal2 s 521078 -960 521190 480 8 la_data_out[112]
port 308 nsew signal output
rlabel metal2 s 524574 -960 524686 480 8 la_data_out[113]
port 309 nsew signal output
rlabel metal2 s 528070 -960 528182 480 8 la_data_out[114]
port 310 nsew signal output
rlabel metal2 s 531658 -960 531770 480 8 la_data_out[115]
port 311 nsew signal output
rlabel metal2 s 535154 -960 535266 480 8 la_data_out[116]
port 312 nsew signal output
rlabel metal2 s 538650 -960 538762 480 8 la_data_out[117]
port 313 nsew signal output
rlabel metal2 s 542238 -960 542350 480 8 la_data_out[118]
port 314 nsew signal output
rlabel metal2 s 545734 -960 545846 480 8 la_data_out[119]
port 315 nsew signal output
rlabel metal2 s 165038 -960 165150 480 8 la_data_out[11]
port 316 nsew signal output
rlabel metal2 s 549230 -960 549342 480 8 la_data_out[120]
port 317 nsew signal output
rlabel metal2 s 552818 -960 552930 480 8 la_data_out[121]
port 318 nsew signal output
rlabel metal2 s 556314 -960 556426 480 8 la_data_out[122]
port 319 nsew signal output
rlabel metal2 s 559810 -960 559922 480 8 la_data_out[123]
port 320 nsew signal output
rlabel metal2 s 563398 -960 563510 480 8 la_data_out[124]
port 321 nsew signal output
rlabel metal2 s 566894 -960 567006 480 8 la_data_out[125]
port 322 nsew signal output
rlabel metal2 s 570390 -960 570502 480 8 la_data_out[126]
port 323 nsew signal output
rlabel metal2 s 573978 -960 574090 480 8 la_data_out[127]
port 324 nsew signal output
rlabel metal2 s 168534 -960 168646 480 8 la_data_out[12]
port 325 nsew signal output
rlabel metal2 s 172030 -960 172142 480 8 la_data_out[13]
port 326 nsew signal output
rlabel metal2 s 175618 -960 175730 480 8 la_data_out[14]
port 327 nsew signal output
rlabel metal2 s 179114 -960 179226 480 8 la_data_out[15]
port 328 nsew signal output
rlabel metal2 s 182610 -960 182722 480 8 la_data_out[16]
port 329 nsew signal output
rlabel metal2 s 186198 -960 186310 480 8 la_data_out[17]
port 330 nsew signal output
rlabel metal2 s 189694 -960 189806 480 8 la_data_out[18]
port 331 nsew signal output
rlabel metal2 s 193190 -960 193302 480 8 la_data_out[19]
port 332 nsew signal output
rlabel metal2 s 129710 -960 129822 480 8 la_data_out[1]
port 333 nsew signal output
rlabel metal2 s 196778 -960 196890 480 8 la_data_out[20]
port 334 nsew signal output
rlabel metal2 s 200274 -960 200386 480 8 la_data_out[21]
port 335 nsew signal output
rlabel metal2 s 203770 -960 203882 480 8 la_data_out[22]
port 336 nsew signal output
rlabel metal2 s 207266 -960 207378 480 8 la_data_out[23]
port 337 nsew signal output
rlabel metal2 s 210854 -960 210966 480 8 la_data_out[24]
port 338 nsew signal output
rlabel metal2 s 214350 -960 214462 480 8 la_data_out[25]
port 339 nsew signal output
rlabel metal2 s 217846 -960 217958 480 8 la_data_out[26]
port 340 nsew signal output
rlabel metal2 s 221434 -960 221546 480 8 la_data_out[27]
port 341 nsew signal output
rlabel metal2 s 224930 -960 225042 480 8 la_data_out[28]
port 342 nsew signal output
rlabel metal2 s 228426 -960 228538 480 8 la_data_out[29]
port 343 nsew signal output
rlabel metal2 s 133298 -960 133410 480 8 la_data_out[2]
port 344 nsew signal output
rlabel metal2 s 232014 -960 232126 480 8 la_data_out[30]
port 345 nsew signal output
rlabel metal2 s 235510 -960 235622 480 8 la_data_out[31]
port 346 nsew signal output
rlabel metal2 s 239006 -960 239118 480 8 la_data_out[32]
port 347 nsew signal output
rlabel metal2 s 242594 -960 242706 480 8 la_data_out[33]
port 348 nsew signal output
rlabel metal2 s 246090 -960 246202 480 8 la_data_out[34]
port 349 nsew signal output
rlabel metal2 s 249586 -960 249698 480 8 la_data_out[35]
port 350 nsew signal output
rlabel metal2 s 253174 -960 253286 480 8 la_data_out[36]
port 351 nsew signal output
rlabel metal2 s 256670 -960 256782 480 8 la_data_out[37]
port 352 nsew signal output
rlabel metal2 s 260166 -960 260278 480 8 la_data_out[38]
port 353 nsew signal output
rlabel metal2 s 263754 -960 263866 480 8 la_data_out[39]
port 354 nsew signal output
rlabel metal2 s 136794 -960 136906 480 8 la_data_out[3]
port 355 nsew signal output
rlabel metal2 s 267250 -960 267362 480 8 la_data_out[40]
port 356 nsew signal output
rlabel metal2 s 270746 -960 270858 480 8 la_data_out[41]
port 357 nsew signal output
rlabel metal2 s 274334 -960 274446 480 8 la_data_out[42]
port 358 nsew signal output
rlabel metal2 s 277830 -960 277942 480 8 la_data_out[43]
port 359 nsew signal output
rlabel metal2 s 281326 -960 281438 480 8 la_data_out[44]
port 360 nsew signal output
rlabel metal2 s 284822 -960 284934 480 8 la_data_out[45]
port 361 nsew signal output
rlabel metal2 s 288410 -960 288522 480 8 la_data_out[46]
port 362 nsew signal output
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[47]
port 363 nsew signal output
rlabel metal2 s 295402 -960 295514 480 8 la_data_out[48]
port 364 nsew signal output
rlabel metal2 s 298990 -960 299102 480 8 la_data_out[49]
port 365 nsew signal output
rlabel metal2 s 140290 -960 140402 480 8 la_data_out[4]
port 366 nsew signal output
rlabel metal2 s 302486 -960 302598 480 8 la_data_out[50]
port 367 nsew signal output
rlabel metal2 s 305982 -960 306094 480 8 la_data_out[51]
port 368 nsew signal output
rlabel metal2 s 309570 -960 309682 480 8 la_data_out[52]
port 369 nsew signal output
rlabel metal2 s 313066 -960 313178 480 8 la_data_out[53]
port 370 nsew signal output
rlabel metal2 s 316562 -960 316674 480 8 la_data_out[54]
port 371 nsew signal output
rlabel metal2 s 320150 -960 320262 480 8 la_data_out[55]
port 372 nsew signal output
rlabel metal2 s 323646 -960 323758 480 8 la_data_out[56]
port 373 nsew signal output
rlabel metal2 s 327142 -960 327254 480 8 la_data_out[57]
port 374 nsew signal output
rlabel metal2 s 330730 -960 330842 480 8 la_data_out[58]
port 375 nsew signal output
rlabel metal2 s 334226 -960 334338 480 8 la_data_out[59]
port 376 nsew signal output
rlabel metal2 s 143878 -960 143990 480 8 la_data_out[5]
port 377 nsew signal output
rlabel metal2 s 337722 -960 337834 480 8 la_data_out[60]
port 378 nsew signal output
rlabel metal2 s 341310 -960 341422 480 8 la_data_out[61]
port 379 nsew signal output
rlabel metal2 s 344806 -960 344918 480 8 la_data_out[62]
port 380 nsew signal output
rlabel metal2 s 348302 -960 348414 480 8 la_data_out[63]
port 381 nsew signal output
rlabel metal2 s 351890 -960 352002 480 8 la_data_out[64]
port 382 nsew signal output
rlabel metal2 s 355386 -960 355498 480 8 la_data_out[65]
port 383 nsew signal output
rlabel metal2 s 358882 -960 358994 480 8 la_data_out[66]
port 384 nsew signal output
rlabel metal2 s 362378 -960 362490 480 8 la_data_out[67]
port 385 nsew signal output
rlabel metal2 s 365966 -960 366078 480 8 la_data_out[68]
port 386 nsew signal output
rlabel metal2 s 369462 -960 369574 480 8 la_data_out[69]
port 387 nsew signal output
rlabel metal2 s 147374 -960 147486 480 8 la_data_out[6]
port 388 nsew signal output
rlabel metal2 s 372958 -960 373070 480 8 la_data_out[70]
port 389 nsew signal output
rlabel metal2 s 376546 -960 376658 480 8 la_data_out[71]
port 390 nsew signal output
rlabel metal2 s 380042 -960 380154 480 8 la_data_out[72]
port 391 nsew signal output
rlabel metal2 s 383538 -960 383650 480 8 la_data_out[73]
port 392 nsew signal output
rlabel metal2 s 387126 -960 387238 480 8 la_data_out[74]
port 393 nsew signal output
rlabel metal2 s 390622 -960 390734 480 8 la_data_out[75]
port 394 nsew signal output
rlabel metal2 s 394118 -960 394230 480 8 la_data_out[76]
port 395 nsew signal output
rlabel metal2 s 397706 -960 397818 480 8 la_data_out[77]
port 396 nsew signal output
rlabel metal2 s 401202 -960 401314 480 8 la_data_out[78]
port 397 nsew signal output
rlabel metal2 s 404698 -960 404810 480 8 la_data_out[79]
port 398 nsew signal output
rlabel metal2 s 150870 -960 150982 480 8 la_data_out[7]
port 399 nsew signal output
rlabel metal2 s 408286 -960 408398 480 8 la_data_out[80]
port 400 nsew signal output
rlabel metal2 s 411782 -960 411894 480 8 la_data_out[81]
port 401 nsew signal output
rlabel metal2 s 415278 -960 415390 480 8 la_data_out[82]
port 402 nsew signal output
rlabel metal2 s 418866 -960 418978 480 8 la_data_out[83]
port 403 nsew signal output
rlabel metal2 s 422362 -960 422474 480 8 la_data_out[84]
port 404 nsew signal output
rlabel metal2 s 425858 -960 425970 480 8 la_data_out[85]
port 405 nsew signal output
rlabel metal2 s 429446 -960 429558 480 8 la_data_out[86]
port 406 nsew signal output
rlabel metal2 s 432942 -960 433054 480 8 la_data_out[87]
port 407 nsew signal output
rlabel metal2 s 436438 -960 436550 480 8 la_data_out[88]
port 408 nsew signal output
rlabel metal2 s 439934 -960 440046 480 8 la_data_out[89]
port 409 nsew signal output
rlabel metal2 s 154458 -960 154570 480 8 la_data_out[8]
port 410 nsew signal output
rlabel metal2 s 443522 -960 443634 480 8 la_data_out[90]
port 411 nsew signal output
rlabel metal2 s 447018 -960 447130 480 8 la_data_out[91]
port 412 nsew signal output
rlabel metal2 s 450514 -960 450626 480 8 la_data_out[92]
port 413 nsew signal output
rlabel metal2 s 454102 -960 454214 480 8 la_data_out[93]
port 414 nsew signal output
rlabel metal2 s 457598 -960 457710 480 8 la_data_out[94]
port 415 nsew signal output
rlabel metal2 s 461094 -960 461206 480 8 la_data_out[95]
port 416 nsew signal output
rlabel metal2 s 464682 -960 464794 480 8 la_data_out[96]
port 417 nsew signal output
rlabel metal2 s 468178 -960 468290 480 8 la_data_out[97]
port 418 nsew signal output
rlabel metal2 s 471674 -960 471786 480 8 la_data_out[98]
port 419 nsew signal output
rlabel metal2 s 475262 -960 475374 480 8 la_data_out[99]
port 420 nsew signal output
rlabel metal2 s 157954 -960 158066 480 8 la_data_out[9]
port 421 nsew signal output
rlabel metal2 s 127410 -960 127522 480 8 la_oen[0]
port 422 nsew signal input
rlabel metal2 s 479954 -960 480066 480 8 la_oen[100]
port 423 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_oen[101]
port 424 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_oen[102]
port 425 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_oen[103]
port 426 nsew signal input
rlabel metal2 s 494030 -960 494142 480 8 la_oen[104]
port 427 nsew signal input
rlabel metal2 s 497526 -960 497638 480 8 la_oen[105]
port 428 nsew signal input
rlabel metal2 s 501114 -960 501226 480 8 la_oen[106]
port 429 nsew signal input
rlabel metal2 s 504610 -960 504722 480 8 la_oen[107]
port 430 nsew signal input
rlabel metal2 s 508106 -960 508218 480 8 la_oen[108]
port 431 nsew signal input
rlabel metal2 s 511694 -960 511806 480 8 la_oen[109]
port 432 nsew signal input
rlabel metal2 s 162646 -960 162758 480 8 la_oen[10]
port 433 nsew signal input
rlabel metal2 s 515190 -960 515302 480 8 la_oen[110]
port 434 nsew signal input
rlabel metal2 s 518686 -960 518798 480 8 la_oen[111]
port 435 nsew signal input
rlabel metal2 s 522274 -960 522386 480 8 la_oen[112]
port 436 nsew signal input
rlabel metal2 s 525770 -960 525882 480 8 la_oen[113]
port 437 nsew signal input
rlabel metal2 s 529266 -960 529378 480 8 la_oen[114]
port 438 nsew signal input
rlabel metal2 s 532854 -960 532966 480 8 la_oen[115]
port 439 nsew signal input
rlabel metal2 s 536350 -960 536462 480 8 la_oen[116]
port 440 nsew signal input
rlabel metal2 s 539846 -960 539958 480 8 la_oen[117]
port 441 nsew signal input
rlabel metal2 s 543342 -960 543454 480 8 la_oen[118]
port 442 nsew signal input
rlabel metal2 s 546930 -960 547042 480 8 la_oen[119]
port 443 nsew signal input
rlabel metal2 s 166142 -960 166254 480 8 la_oen[11]
port 444 nsew signal input
rlabel metal2 s 550426 -960 550538 480 8 la_oen[120]
port 445 nsew signal input
rlabel metal2 s 553922 -960 554034 480 8 la_oen[121]
port 446 nsew signal input
rlabel metal2 s 557510 -960 557622 480 8 la_oen[122]
port 447 nsew signal input
rlabel metal2 s 561006 -960 561118 480 8 la_oen[123]
port 448 nsew signal input
rlabel metal2 s 564502 -960 564614 480 8 la_oen[124]
port 449 nsew signal input
rlabel metal2 s 568090 -960 568202 480 8 la_oen[125]
port 450 nsew signal input
rlabel metal2 s 571586 -960 571698 480 8 la_oen[126]
port 451 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oen[127]
port 452 nsew signal input
rlabel metal2 s 169730 -960 169842 480 8 la_oen[12]
port 453 nsew signal input
rlabel metal2 s 173226 -960 173338 480 8 la_oen[13]
port 454 nsew signal input
rlabel metal2 s 176722 -960 176834 480 8 la_oen[14]
port 455 nsew signal input
rlabel metal2 s 180310 -960 180422 480 8 la_oen[15]
port 456 nsew signal input
rlabel metal2 s 183806 -960 183918 480 8 la_oen[16]
port 457 nsew signal input
rlabel metal2 s 187302 -960 187414 480 8 la_oen[17]
port 458 nsew signal input
rlabel metal2 s 190890 -960 191002 480 8 la_oen[18]
port 459 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_oen[19]
port 460 nsew signal input
rlabel metal2 s 130906 -960 131018 480 8 la_oen[1]
port 461 nsew signal input
rlabel metal2 s 197882 -960 197994 480 8 la_oen[20]
port 462 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_oen[21]
port 463 nsew signal input
rlabel metal2 s 204966 -960 205078 480 8 la_oen[22]
port 464 nsew signal input
rlabel metal2 s 208462 -960 208574 480 8 la_oen[23]
port 465 nsew signal input
rlabel metal2 s 212050 -960 212162 480 8 la_oen[24]
port 466 nsew signal input
rlabel metal2 s 215546 -960 215658 480 8 la_oen[25]
port 467 nsew signal input
rlabel metal2 s 219042 -960 219154 480 8 la_oen[26]
port 468 nsew signal input
rlabel metal2 s 222630 -960 222742 480 8 la_oen[27]
port 469 nsew signal input
rlabel metal2 s 226126 -960 226238 480 8 la_oen[28]
port 470 nsew signal input
rlabel metal2 s 229622 -960 229734 480 8 la_oen[29]
port 471 nsew signal input
rlabel metal2 s 134494 -960 134606 480 8 la_oen[2]
port 472 nsew signal input
rlabel metal2 s 233118 -960 233230 480 8 la_oen[30]
port 473 nsew signal input
rlabel metal2 s 236706 -960 236818 480 8 la_oen[31]
port 474 nsew signal input
rlabel metal2 s 240202 -960 240314 480 8 la_oen[32]
port 475 nsew signal input
rlabel metal2 s 243698 -960 243810 480 8 la_oen[33]
port 476 nsew signal input
rlabel metal2 s 247286 -960 247398 480 8 la_oen[34]
port 477 nsew signal input
rlabel metal2 s 250782 -960 250894 480 8 la_oen[35]
port 478 nsew signal input
rlabel metal2 s 254278 -960 254390 480 8 la_oen[36]
port 479 nsew signal input
rlabel metal2 s 257866 -960 257978 480 8 la_oen[37]
port 480 nsew signal input
rlabel metal2 s 261362 -960 261474 480 8 la_oen[38]
port 481 nsew signal input
rlabel metal2 s 264858 -960 264970 480 8 la_oen[39]
port 482 nsew signal input
rlabel metal2 s 137990 -960 138102 480 8 la_oen[3]
port 483 nsew signal input
rlabel metal2 s 268446 -960 268558 480 8 la_oen[40]
port 484 nsew signal input
rlabel metal2 s 271942 -960 272054 480 8 la_oen[41]
port 485 nsew signal input
rlabel metal2 s 275438 -960 275550 480 8 la_oen[42]
port 486 nsew signal input
rlabel metal2 s 279026 -960 279138 480 8 la_oen[43]
port 487 nsew signal input
rlabel metal2 s 282522 -960 282634 480 8 la_oen[44]
port 488 nsew signal input
rlabel metal2 s 286018 -960 286130 480 8 la_oen[45]
port 489 nsew signal input
rlabel metal2 s 289606 -960 289718 480 8 la_oen[46]
port 490 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[47]
port 491 nsew signal input
rlabel metal2 s 296598 -960 296710 480 8 la_oen[48]
port 492 nsew signal input
rlabel metal2 s 300186 -960 300298 480 8 la_oen[49]
port 493 nsew signal input
rlabel metal2 s 141486 -960 141598 480 8 la_oen[4]
port 494 nsew signal input
rlabel metal2 s 303682 -960 303794 480 8 la_oen[50]
port 495 nsew signal input
rlabel metal2 s 307178 -960 307290 480 8 la_oen[51]
port 496 nsew signal input
rlabel metal2 s 310674 -960 310786 480 8 la_oen[52]
port 497 nsew signal input
rlabel metal2 s 314262 -960 314374 480 8 la_oen[53]
port 498 nsew signal input
rlabel metal2 s 317758 -960 317870 480 8 la_oen[54]
port 499 nsew signal input
rlabel metal2 s 321254 -960 321366 480 8 la_oen[55]
port 500 nsew signal input
rlabel metal2 s 324842 -960 324954 480 8 la_oen[56]
port 501 nsew signal input
rlabel metal2 s 328338 -960 328450 480 8 la_oen[57]
port 502 nsew signal input
rlabel metal2 s 331834 -960 331946 480 8 la_oen[58]
port 503 nsew signal input
rlabel metal2 s 335422 -960 335534 480 8 la_oen[59]
port 504 nsew signal input
rlabel metal2 s 145074 -960 145186 480 8 la_oen[5]
port 505 nsew signal input
rlabel metal2 s 338918 -960 339030 480 8 la_oen[60]
port 506 nsew signal input
rlabel metal2 s 342414 -960 342526 480 8 la_oen[61]
port 507 nsew signal input
rlabel metal2 s 346002 -960 346114 480 8 la_oen[62]
port 508 nsew signal input
rlabel metal2 s 349498 -960 349610 480 8 la_oen[63]
port 509 nsew signal input
rlabel metal2 s 352994 -960 353106 480 8 la_oen[64]
port 510 nsew signal input
rlabel metal2 s 356582 -960 356694 480 8 la_oen[65]
port 511 nsew signal input
rlabel metal2 s 360078 -960 360190 480 8 la_oen[66]
port 512 nsew signal input
rlabel metal2 s 363574 -960 363686 480 8 la_oen[67]
port 513 nsew signal input
rlabel metal2 s 367162 -960 367274 480 8 la_oen[68]
port 514 nsew signal input
rlabel metal2 s 370658 -960 370770 480 8 la_oen[69]
port 515 nsew signal input
rlabel metal2 s 148570 -960 148682 480 8 la_oen[6]
port 516 nsew signal input
rlabel metal2 s 374154 -960 374266 480 8 la_oen[70]
port 517 nsew signal input
rlabel metal2 s 377742 -960 377854 480 8 la_oen[71]
port 518 nsew signal input
rlabel metal2 s 381238 -960 381350 480 8 la_oen[72]
port 519 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_oen[73]
port 520 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_oen[74]
port 521 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_oen[75]
port 522 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_oen[76]
port 523 nsew signal input
rlabel metal2 s 398810 -960 398922 480 8 la_oen[77]
port 524 nsew signal input
rlabel metal2 s 402398 -960 402510 480 8 la_oen[78]
port 525 nsew signal input
rlabel metal2 s 405894 -960 406006 480 8 la_oen[79]
port 526 nsew signal input
rlabel metal2 s 152066 -960 152178 480 8 la_oen[7]
port 527 nsew signal input
rlabel metal2 s 409390 -960 409502 480 8 la_oen[80]
port 528 nsew signal input
rlabel metal2 s 412978 -960 413090 480 8 la_oen[81]
port 529 nsew signal input
rlabel metal2 s 416474 -960 416586 480 8 la_oen[82]
port 530 nsew signal input
rlabel metal2 s 419970 -960 420082 480 8 la_oen[83]
port 531 nsew signal input
rlabel metal2 s 423558 -960 423670 480 8 la_oen[84]
port 532 nsew signal input
rlabel metal2 s 427054 -960 427166 480 8 la_oen[85]
port 533 nsew signal input
rlabel metal2 s 430550 -960 430662 480 8 la_oen[86]
port 534 nsew signal input
rlabel metal2 s 434138 -960 434250 480 8 la_oen[87]
port 535 nsew signal input
rlabel metal2 s 437634 -960 437746 480 8 la_oen[88]
port 536 nsew signal input
rlabel metal2 s 441130 -960 441242 480 8 la_oen[89]
port 537 nsew signal input
rlabel metal2 s 155562 -960 155674 480 8 la_oen[8]
port 538 nsew signal input
rlabel metal2 s 444718 -960 444830 480 8 la_oen[90]
port 539 nsew signal input
rlabel metal2 s 448214 -960 448326 480 8 la_oen[91]
port 540 nsew signal input
rlabel metal2 s 451710 -960 451822 480 8 la_oen[92]
port 541 nsew signal input
rlabel metal2 s 455298 -960 455410 480 8 la_oen[93]
port 542 nsew signal input
rlabel metal2 s 458794 -960 458906 480 8 la_oen[94]
port 543 nsew signal input
rlabel metal2 s 462290 -960 462402 480 8 la_oen[95]
port 544 nsew signal input
rlabel metal2 s 465786 -960 465898 480 8 la_oen[96]
port 545 nsew signal input
rlabel metal2 s 469374 -960 469486 480 8 la_oen[97]
port 546 nsew signal input
rlabel metal2 s 472870 -960 472982 480 8 la_oen[98]
port 547 nsew signal input
rlabel metal2 s 476366 -960 476478 480 8 la_oen[99]
port 548 nsew signal input
rlabel metal2 s 159150 -960 159262 480 8 la_oen[9]
port 549 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 user_clock2
port 550 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 551 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 552 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 553 nsew signal output
rlabel metal2 s 7534 -960 7646 480 8 wbs_adr_i[0]
port 554 nsew signal input
rlabel metal2 s 47462 -960 47574 480 8 wbs_adr_i[10]
port 555 nsew signal input
rlabel metal2 s 51050 -960 51162 480 8 wbs_adr_i[11]
port 556 nsew signal input
rlabel metal2 s 54546 -960 54658 480 8 wbs_adr_i[12]
port 557 nsew signal input
rlabel metal2 s 58042 -960 58154 480 8 wbs_adr_i[13]
port 558 nsew signal input
rlabel metal2 s 61630 -960 61742 480 8 wbs_adr_i[14]
port 559 nsew signal input
rlabel metal2 s 65126 -960 65238 480 8 wbs_adr_i[15]
port 560 nsew signal input
rlabel metal2 s 68622 -960 68734 480 8 wbs_adr_i[16]
port 561 nsew signal input
rlabel metal2 s 72210 -960 72322 480 8 wbs_adr_i[17]
port 562 nsew signal input
rlabel metal2 s 75706 -960 75818 480 8 wbs_adr_i[18]
port 563 nsew signal input
rlabel metal2 s 79202 -960 79314 480 8 wbs_adr_i[19]
port 564 nsew signal input
rlabel metal2 s 12226 -960 12338 480 8 wbs_adr_i[1]
port 565 nsew signal input
rlabel metal2 s 82790 -960 82902 480 8 wbs_adr_i[20]
port 566 nsew signal input
rlabel metal2 s 86286 -960 86398 480 8 wbs_adr_i[21]
port 567 nsew signal input
rlabel metal2 s 89782 -960 89894 480 8 wbs_adr_i[22]
port 568 nsew signal input
rlabel metal2 s 93370 -960 93482 480 8 wbs_adr_i[23]
port 569 nsew signal input
rlabel metal2 s 96866 -960 96978 480 8 wbs_adr_i[24]
port 570 nsew signal input
rlabel metal2 s 100362 -960 100474 480 8 wbs_adr_i[25]
port 571 nsew signal input
rlabel metal2 s 103858 -960 103970 480 8 wbs_adr_i[26]
port 572 nsew signal input
rlabel metal2 s 107446 -960 107558 480 8 wbs_adr_i[27]
port 573 nsew signal input
rlabel metal2 s 110942 -960 111054 480 8 wbs_adr_i[28]
port 574 nsew signal input
rlabel metal2 s 114438 -960 114550 480 8 wbs_adr_i[29]
port 575 nsew signal input
rlabel metal2 s 16918 -960 17030 480 8 wbs_adr_i[2]
port 576 nsew signal input
rlabel metal2 s 118026 -960 118138 480 8 wbs_adr_i[30]
port 577 nsew signal input
rlabel metal2 s 121522 -960 121634 480 8 wbs_adr_i[31]
port 578 nsew signal input
rlabel metal2 s 21610 -960 21722 480 8 wbs_adr_i[3]
port 579 nsew signal input
rlabel metal2 s 26302 -960 26414 480 8 wbs_adr_i[4]
port 580 nsew signal input
rlabel metal2 s 29890 -960 30002 480 8 wbs_adr_i[5]
port 581 nsew signal input
rlabel metal2 s 33386 -960 33498 480 8 wbs_adr_i[6]
port 582 nsew signal input
rlabel metal2 s 36882 -960 36994 480 8 wbs_adr_i[7]
port 583 nsew signal input
rlabel metal2 s 40470 -960 40582 480 8 wbs_adr_i[8]
port 584 nsew signal input
rlabel metal2 s 43966 -960 44078 480 8 wbs_adr_i[9]
port 585 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 586 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 587 nsew signal input
rlabel metal2 s 48658 -960 48770 480 8 wbs_dat_i[10]
port 588 nsew signal input
rlabel metal2 s 52154 -960 52266 480 8 wbs_dat_i[11]
port 589 nsew signal input
rlabel metal2 s 55742 -960 55854 480 8 wbs_dat_i[12]
port 590 nsew signal input
rlabel metal2 s 59238 -960 59350 480 8 wbs_dat_i[13]
port 591 nsew signal input
rlabel metal2 s 62734 -960 62846 480 8 wbs_dat_i[14]
port 592 nsew signal input
rlabel metal2 s 66322 -960 66434 480 8 wbs_dat_i[15]
port 593 nsew signal input
rlabel metal2 s 69818 -960 69930 480 8 wbs_dat_i[16]
port 594 nsew signal input
rlabel metal2 s 73314 -960 73426 480 8 wbs_dat_i[17]
port 595 nsew signal input
rlabel metal2 s 76902 -960 77014 480 8 wbs_dat_i[18]
port 596 nsew signal input
rlabel metal2 s 80398 -960 80510 480 8 wbs_dat_i[19]
port 597 nsew signal input
rlabel metal2 s 13422 -960 13534 480 8 wbs_dat_i[1]
port 598 nsew signal input
rlabel metal2 s 83894 -960 84006 480 8 wbs_dat_i[20]
port 599 nsew signal input
rlabel metal2 s 87482 -960 87594 480 8 wbs_dat_i[21]
port 600 nsew signal input
rlabel metal2 s 90978 -960 91090 480 8 wbs_dat_i[22]
port 601 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_dat_i[23]
port 602 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_dat_i[24]
port 603 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_dat_i[25]
port 604 nsew signal input
rlabel metal2 s 105054 -960 105166 480 8 wbs_dat_i[26]
port 605 nsew signal input
rlabel metal2 s 108642 -960 108754 480 8 wbs_dat_i[27]
port 606 nsew signal input
rlabel metal2 s 112138 -960 112250 480 8 wbs_dat_i[28]
port 607 nsew signal input
rlabel metal2 s 115634 -960 115746 480 8 wbs_dat_i[29]
port 608 nsew signal input
rlabel metal2 s 18114 -960 18226 480 8 wbs_dat_i[2]
port 609 nsew signal input
rlabel metal2 s 119222 -960 119334 480 8 wbs_dat_i[30]
port 610 nsew signal input
rlabel metal2 s 122718 -960 122830 480 8 wbs_dat_i[31]
port 611 nsew signal input
rlabel metal2 s 22806 -960 22918 480 8 wbs_dat_i[3]
port 612 nsew signal input
rlabel metal2 s 27498 -960 27610 480 8 wbs_dat_i[4]
port 613 nsew signal input
rlabel metal2 s 31086 -960 31198 480 8 wbs_dat_i[5]
port 614 nsew signal input
rlabel metal2 s 34582 -960 34694 480 8 wbs_dat_i[6]
port 615 nsew signal input
rlabel metal2 s 38078 -960 38190 480 8 wbs_dat_i[7]
port 616 nsew signal input
rlabel metal2 s 41666 -960 41778 480 8 wbs_dat_i[8]
port 617 nsew signal input
rlabel metal2 s 45162 -960 45274 480 8 wbs_dat_i[9]
port 618 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 619 nsew signal output
rlabel metal2 s 49854 -960 49966 480 8 wbs_dat_o[10]
port 620 nsew signal output
rlabel metal2 s 53350 -960 53462 480 8 wbs_dat_o[11]
port 621 nsew signal output
rlabel metal2 s 56938 -960 57050 480 8 wbs_dat_o[12]
port 622 nsew signal output
rlabel metal2 s 60434 -960 60546 480 8 wbs_dat_o[13]
port 623 nsew signal output
rlabel metal2 s 63930 -960 64042 480 8 wbs_dat_o[14]
port 624 nsew signal output
rlabel metal2 s 67518 -960 67630 480 8 wbs_dat_o[15]
port 625 nsew signal output
rlabel metal2 s 71014 -960 71126 480 8 wbs_dat_o[16]
port 626 nsew signal output
rlabel metal2 s 74510 -960 74622 480 8 wbs_dat_o[17]
port 627 nsew signal output
rlabel metal2 s 78006 -960 78118 480 8 wbs_dat_o[18]
port 628 nsew signal output
rlabel metal2 s 81594 -960 81706 480 8 wbs_dat_o[19]
port 629 nsew signal output
rlabel metal2 s 14618 -960 14730 480 8 wbs_dat_o[1]
port 630 nsew signal output
rlabel metal2 s 85090 -960 85202 480 8 wbs_dat_o[20]
port 631 nsew signal output
rlabel metal2 s 88586 -960 88698 480 8 wbs_dat_o[21]
port 632 nsew signal output
rlabel metal2 s 92174 -960 92286 480 8 wbs_dat_o[22]
port 633 nsew signal output
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_o[23]
port 634 nsew signal output
rlabel metal2 s 99166 -960 99278 480 8 wbs_dat_o[24]
port 635 nsew signal output
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_o[25]
port 636 nsew signal output
rlabel metal2 s 106250 -960 106362 480 8 wbs_dat_o[26]
port 637 nsew signal output
rlabel metal2 s 109746 -960 109858 480 8 wbs_dat_o[27]
port 638 nsew signal output
rlabel metal2 s 113334 -960 113446 480 8 wbs_dat_o[28]
port 639 nsew signal output
rlabel metal2 s 116830 -960 116942 480 8 wbs_dat_o[29]
port 640 nsew signal output
rlabel metal2 s 19310 -960 19422 480 8 wbs_dat_o[2]
port 641 nsew signal output
rlabel metal2 s 120326 -960 120438 480 8 wbs_dat_o[30]
port 642 nsew signal output
rlabel metal2 s 123914 -960 124026 480 8 wbs_dat_o[31]
port 643 nsew signal output
rlabel metal2 s 24002 -960 24114 480 8 wbs_dat_o[3]
port 644 nsew signal output
rlabel metal2 s 28694 -960 28806 480 8 wbs_dat_o[4]
port 645 nsew signal output
rlabel metal2 s 32190 -960 32302 480 8 wbs_dat_o[5]
port 646 nsew signal output
rlabel metal2 s 35778 -960 35890 480 8 wbs_dat_o[6]
port 647 nsew signal output
rlabel metal2 s 39274 -960 39386 480 8 wbs_dat_o[7]
port 648 nsew signal output
rlabel metal2 s 42770 -960 42882 480 8 wbs_dat_o[8]
port 649 nsew signal output
rlabel metal2 s 46358 -960 46470 480 8 wbs_dat_o[9]
port 650 nsew signal output
rlabel metal2 s 11030 -960 11142 480 8 wbs_sel_i[0]
port 651 nsew signal input
rlabel metal2 s 15814 -960 15926 480 8 wbs_sel_i[1]
port 652 nsew signal input
rlabel metal2 s 20506 -960 20618 480 8 wbs_sel_i[2]
port 653 nsew signal input
rlabel metal2 s 25198 -960 25310 480 8 wbs_sel_i[3]
port 654 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 655 nsew signal input
rlabel metal2 s 6338 -960 6450 480 8 wbs_we_i
port 656 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 705800 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 705800 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 705800 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 705800 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 705800 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 705800 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 325804 459952 326404 705800 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 289804 459952 290404 705800 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 253804 459952 254404 705800 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 705800 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 705800 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 705800 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 705800 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 705800 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 705800 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 336048 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 336048 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 336048 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s -2936 686828 586860 687428 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s -2936 650828 586860 651428 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s -2936 614828 586860 615428 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s -2936 578828 586860 579428 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s -2936 542828 586860 543428 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s -2936 506828 586860 507428 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s -2936 470828 586860 471428 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s -2936 434828 586860 435428 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s -2936 398828 586860 399428 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s -2936 362828 586860 363428 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s -2936 326828 586860 327428 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s -2936 290828 586860 291428 6 vccd1
port 691 nsew power bidirectional
rlabel metal5 s -2936 254828 586860 255428 6 vccd1
port 692 nsew power bidirectional
rlabel metal5 s -2936 218828 586860 219428 6 vccd1
port 693 nsew power bidirectional
rlabel metal5 s -2936 182828 586860 183428 6 vccd1
port 694 nsew power bidirectional
rlabel metal5 s -2936 146828 586860 147428 6 vccd1
port 695 nsew power bidirectional
rlabel metal5 s -2936 110828 586860 111428 6 vccd1
port 696 nsew power bidirectional
rlabel metal5 s -2936 74828 586860 75428 6 vccd1
port 697 nsew power bidirectional
rlabel metal5 s -2936 38828 586860 39428 6 vccd1
port 698 nsew power bidirectional
rlabel metal5 s -2936 2828 586860 3428 6 vccd1
port 699 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 700 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 705800 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 705800 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 705800 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 705800 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 705800 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 705800 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 343804 459952 344404 705800 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 307804 459952 308404 705800 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s 271804 459952 272404 705800 6 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 235804 459952 236404 705800 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 705800 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 705800 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 705800 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 705800 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 705800 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 705800 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 336048 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 336048 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 336048 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 336048 6 vssd1
port 722 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 723 nsew ground bidirectional
rlabel metal5 s -2936 668828 586860 669428 6 vssd1
port 724 nsew ground bidirectional
rlabel metal5 s -2936 632828 586860 633428 6 vssd1
port 725 nsew ground bidirectional
rlabel metal5 s -2936 596828 586860 597428 6 vssd1
port 726 nsew ground bidirectional
rlabel metal5 s -2936 560828 586860 561428 6 vssd1
port 727 nsew ground bidirectional
rlabel metal5 s -2936 524828 586860 525428 6 vssd1
port 728 nsew ground bidirectional
rlabel metal5 s -2936 488828 586860 489428 6 vssd1
port 729 nsew ground bidirectional
rlabel metal5 s -2936 452828 586860 453428 6 vssd1
port 730 nsew ground bidirectional
rlabel metal5 s -2936 416828 586860 417428 6 vssd1
port 731 nsew ground bidirectional
rlabel metal5 s -2936 380828 586860 381428 6 vssd1
port 732 nsew ground bidirectional
rlabel metal5 s -2936 344828 586860 345428 6 vssd1
port 733 nsew ground bidirectional
rlabel metal5 s -2936 308828 586860 309428 6 vssd1
port 734 nsew ground bidirectional
rlabel metal5 s -2936 272828 586860 273428 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s -2936 236828 586860 237428 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s -2936 200828 586860 201428 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s -2936 164828 586860 165428 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s -2936 128828 586860 129428 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s -2936 92828 586860 93428 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s -2936 56828 586860 57428 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s -2936 20828 586860 21428 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 744 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 707680 6 vccd2
port 745 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 707680 6 vccd2
port 746 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 707680 6 vccd2
port 747 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 707680 6 vccd2
port 748 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 707680 6 vccd2
port 749 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 707680 6 vccd2
port 750 nsew power bidirectional
rlabel metal4 s 329404 460000 330004 707680 6 vccd2
port 751 nsew power bidirectional
rlabel metal4 s 293404 460000 294004 707680 6 vccd2
port 752 nsew power bidirectional
rlabel metal4 s 257404 460000 258004 707680 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 707680 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 707680 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 707680 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 707680 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 707680 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 707680 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 336000 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 336000 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 336000 6 vccd2
port 765 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 766 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 767 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 768 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 769 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 770 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 771 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 772 nsew power bidirectional
rlabel metal5 s -4816 474476 588740 475076 6 vccd2
port 773 nsew power bidirectional
rlabel metal5 s -4816 438476 588740 439076 6 vccd2
port 774 nsew power bidirectional
rlabel metal5 s -4816 402476 588740 403076 6 vccd2
port 775 nsew power bidirectional
rlabel metal5 s -4816 366476 588740 367076 6 vccd2
port 776 nsew power bidirectional
rlabel metal5 s -4816 330476 588740 331076 6 vccd2
port 777 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 778 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 779 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 780 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 781 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 782 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 783 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 784 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 785 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 786 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 787 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 788 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 707680 6 vssd2
port 789 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 707680 6 vssd2
port 790 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 707680 6 vssd2
port 791 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 707680 6 vssd2
port 792 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 707680 6 vssd2
port 793 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 707680 6 vssd2
port 794 nsew ground bidirectional
rlabel metal4 s 347404 460000 348004 707680 6 vssd2
port 795 nsew ground bidirectional
rlabel metal4 s 311404 460000 312004 707680 6 vssd2
port 796 nsew ground bidirectional
rlabel metal4 s 275404 460000 276004 707680 6 vssd2
port 797 nsew ground bidirectional
rlabel metal4 s 239404 460000 240004 707680 6 vssd2
port 798 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 707680 6 vssd2
port 799 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 707680 6 vssd2
port 800 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 707680 6 vssd2
port 801 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 707680 6 vssd2
port 802 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 707680 6 vssd2
port 803 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 336000 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 336000 6 vssd2
port 807 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 336000 6 vssd2
port 808 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 336000 6 vssd2
port 809 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 810 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 811 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 812 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 813 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 814 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 815 nsew ground bidirectional
rlabel metal5 s -4816 492476 588740 493076 6 vssd2
port 816 nsew ground bidirectional
rlabel metal5 s -4816 456476 588740 457076 6 vssd2
port 817 nsew ground bidirectional
rlabel metal5 s -4816 420476 588740 421076 6 vssd2
port 818 nsew ground bidirectional
rlabel metal5 s -4816 384476 588740 385076 6 vssd2
port 819 nsew ground bidirectional
rlabel metal5 s -4816 348476 588740 349076 6 vssd2
port 820 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 821 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 822 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 823 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 824 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 825 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 826 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 827 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 828 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 829 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 830 nsew ground bidirectional
rlabel metal4 s 549004 -5624 549604 709560 6 vdda1
port 831 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 709560 6 vdda1
port 832 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 709560 6 vdda1
port 833 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 709560 6 vdda1
port 834 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 709560 6 vdda1
port 835 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 709560 6 vdda1
port 836 nsew power bidirectional
rlabel metal4 s 333004 460000 333604 709560 6 vdda1
port 837 nsew power bidirectional
rlabel metal4 s 297004 460000 297604 709560 6 vdda1
port 838 nsew power bidirectional
rlabel metal4 s 261004 460000 261604 709560 6 vdda1
port 839 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 709560 6 vdda1
port 840 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 709560 6 vdda1
port 841 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 709560 6 vdda1
port 842 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 709560 6 vdda1
port 843 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 709560 6 vdda1
port 844 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 709560 6 vdda1
port 845 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 846 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 847 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 848 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 336000 6 vdda1
port 849 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 336000 6 vdda1
port 850 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 336000 6 vdda1
port 851 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 852 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 853 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 854 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 855 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 856 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 857 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 858 nsew power bidirectional
rlabel metal5 s -6696 478076 590620 478676 6 vdda1
port 859 nsew power bidirectional
rlabel metal5 s -6696 442076 590620 442676 6 vdda1
port 860 nsew power bidirectional
rlabel metal5 s -6696 406076 590620 406676 6 vdda1
port 861 nsew power bidirectional
rlabel metal5 s -6696 370076 590620 370676 6 vdda1
port 862 nsew power bidirectional
rlabel metal5 s -6696 334076 590620 334676 6 vdda1
port 863 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 864 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 865 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 866 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 867 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 868 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 869 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 870 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 871 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 872 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 873 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 874 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1
port 875 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 709560 6 vssa1
port 876 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 709560 6 vssa1
port 877 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 709560 6 vssa1
port 878 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 709560 6 vssa1
port 879 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 709560 6 vssa1
port 880 nsew ground bidirectional
rlabel metal4 s 351004 460000 351604 709560 6 vssa1
port 881 nsew ground bidirectional
rlabel metal4 s 315004 460000 315604 709560 6 vssa1
port 882 nsew ground bidirectional
rlabel metal4 s 279004 460000 279604 709560 6 vssa1
port 883 nsew ground bidirectional
rlabel metal4 s 243004 460000 243604 709560 6 vssa1
port 884 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 709560 6 vssa1
port 885 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 709560 6 vssa1
port 886 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 709560 6 vssa1
port 887 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 709560 6 vssa1
port 888 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 709560 6 vssa1
port 889 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1
port 890 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 891 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 336000 6 vssa1
port 892 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 336000 6 vssa1
port 893 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 336000 6 vssa1
port 894 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 336000 6 vssa1
port 895 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 896 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 897 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 898 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 899 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 900 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 901 nsew ground bidirectional
rlabel metal5 s -6696 496076 590620 496676 6 vssa1
port 902 nsew ground bidirectional
rlabel metal5 s -6696 460076 590620 460676 6 vssa1
port 903 nsew ground bidirectional
rlabel metal5 s -6696 424076 590620 424676 6 vssa1
port 904 nsew ground bidirectional
rlabel metal5 s -6696 388076 590620 388676 6 vssa1
port 905 nsew ground bidirectional
rlabel metal5 s -6696 352076 590620 352676 6 vssa1
port 906 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 907 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 908 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 909 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 910 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 911 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 912 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 913 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 914 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 915 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 916 nsew ground bidirectional
rlabel metal4 s 552604 -7504 553204 711440 6 vdda2
port 917 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 711440 6 vdda2
port 918 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 711440 6 vdda2
port 919 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 711440 6 vdda2
port 920 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 711440 6 vdda2
port 921 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 711440 6 vdda2
port 922 nsew power bidirectional
rlabel metal4 s 336604 460000 337204 711440 6 vdda2
port 923 nsew power bidirectional
rlabel metal4 s 300604 460000 301204 711440 6 vdda2
port 924 nsew power bidirectional
rlabel metal4 s 264604 460000 265204 711440 6 vdda2
port 925 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 711440 6 vdda2
port 926 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 711440 6 vdda2
port 927 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 711440 6 vdda2
port 928 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 711440 6 vdda2
port 929 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 711440 6 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 711440 6 vdda2
port 931 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 932 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 933 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 934 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 336000 6 vdda2
port 935 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 336000 6 vdda2
port 936 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 336000 6 vdda2
port 937 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 938 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 939 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 940 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 941 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 942 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 943 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 944 nsew power bidirectional
rlabel metal5 s -8576 481676 592500 482276 6 vdda2
port 945 nsew power bidirectional
rlabel metal5 s -8576 445676 592500 446276 6 vdda2
port 946 nsew power bidirectional
rlabel metal5 s -8576 409676 592500 410276 6 vdda2
port 947 nsew power bidirectional
rlabel metal5 s -8576 373676 592500 374276 6 vdda2
port 948 nsew power bidirectional
rlabel metal5 s -8576 337676 592500 338276 6 vdda2
port 949 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 950 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 951 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 952 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 953 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 954 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 955 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 956 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 957 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 958 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 959 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 960 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2
port 961 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 711440 6 vssa2
port 962 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 711440 6 vssa2
port 963 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 711440 6 vssa2
port 964 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 711440 6 vssa2
port 965 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 711440 6 vssa2
port 966 nsew ground bidirectional
rlabel metal4 s 354604 460000 355204 711440 6 vssa2
port 967 nsew ground bidirectional
rlabel metal4 s 318604 460000 319204 711440 6 vssa2
port 968 nsew ground bidirectional
rlabel metal4 s 282604 460000 283204 711440 6 vssa2
port 969 nsew ground bidirectional
rlabel metal4 s 246604 460000 247204 711440 6 vssa2
port 970 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 711440 6 vssa2
port 971 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 711440 6 vssa2
port 972 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 711440 6 vssa2
port 973 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 711440 6 vssa2
port 974 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 711440 6 vssa2
port 975 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2
port 976 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 977 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 336000 6 vssa2
port 978 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 336000 6 vssa2
port 979 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 336000 6 vssa2
port 980 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 336000 6 vssa2
port 981 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 982 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 983 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 984 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 985 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 986 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 987 nsew ground bidirectional
rlabel metal5 s -8576 499676 592500 500276 6 vssa2
port 988 nsew ground bidirectional
rlabel metal5 s -8576 463676 592500 464276 6 vssa2
port 989 nsew ground bidirectional
rlabel metal5 s -8576 427676 592500 428276 6 vssa2
port 990 nsew ground bidirectional
rlabel metal5 s -8576 391676 592500 392276 6 vssa2
port 991 nsew ground bidirectional
rlabel metal5 s -8576 355676 592500 356276 6 vssa2
port 992 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 993 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 994 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 995 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 996 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 997 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 998 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 999 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 1000 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 1001 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1002 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 40990274
string GDS_START 6085648
<< end >>

