magic
tech sky130A
magscale 1 2
timestamp 1640931048
<< nwell >>
rect 0 11 974 384
rect 1153 11 1742 384
<< pwell >>
rect 184 474 763 848
rect 966 452 1811 958
<< locali >>
rect 569 379 655 417
rect 591 363 655 379
rect 592 330 655 363
rect 592 327 668 330
rect 592 310 713 327
rect 592 276 662 310
rect 696 276 713 310
rect 592 265 713 276
rect 592 264 668 265
<< viali >>
rect 2196 852 2230 886
rect 357 381 391 415
rect 1624 406 1658 440
rect 1838 412 1872 446
rect 2098 310 2132 344
rect 662 276 696 310
rect 172 204 206 238
<< metal1 >>
rect -1 1331 243 1430
rect 644 894 718 900
rect 2186 894 2242 900
rect 644 840 650 894
rect 712 886 2242 894
rect 712 852 2196 886
rect 2230 852 2242 886
rect 712 842 2242 852
rect 712 840 718 842
rect 644 834 718 840
rect 2186 838 2242 842
rect 66 458 130 464
rect 66 404 72 458
rect 124 404 130 458
rect 1474 440 1674 458
rect 2180 456 2246 462
rect 2180 454 2186 456
rect 66 398 130 404
rect 338 415 416 416
rect 338 381 357 415
rect 391 381 416 415
rect 1474 406 1624 440
rect 1658 406 1674 440
rect 1474 390 1674 406
rect 1826 446 2186 454
rect 1826 412 1838 446
rect 1872 412 2186 446
rect 1826 404 2186 412
rect 2240 404 2246 456
rect 2180 398 2246 404
rect 338 366 416 381
rect 2084 344 2300 354
rect 648 324 712 330
rect 648 270 654 324
rect 706 270 712 324
rect 2084 310 2098 344
rect 2132 310 2300 344
rect 2084 302 2300 310
rect 648 264 712 270
rect 64 250 128 252
rect 64 246 216 250
rect 64 194 70 246
rect 122 238 216 246
rect 122 204 172 238
rect 206 204 216 238
rect 122 194 216 204
rect 64 190 216 194
rect 64 188 128 190
rect 11 74 828 98
rect 11 24 846 74
rect 11 0 836 24
rect 1478 0 1594 98
<< via1 >>
rect 650 840 712 894
rect 72 404 124 458
rect 2186 404 2240 456
rect 654 310 706 324
rect 654 276 662 310
rect 662 276 696 310
rect 696 276 706 310
rect 654 270 706 276
rect 70 194 122 246
<< metal2 >>
rect 68 464 128 1434
rect 2184 1020 2238 1430
rect 644 894 718 900
rect 644 840 650 894
rect 712 840 718 894
rect 644 834 718 840
rect 66 458 130 464
rect 66 404 72 458
rect 124 404 130 458
rect 66 398 130 404
rect 650 330 710 834
rect 2180 456 2246 462
rect 2180 404 2186 456
rect 2240 404 2246 456
rect 2180 398 2246 404
rect 648 324 712 330
rect 648 270 654 324
rect 706 270 712 324
rect 648 264 712 270
rect 64 246 128 252
rect 64 194 70 246
rect 122 194 128 246
rect 64 188 128 194
rect 68 0 128 188
rect 2184 0 2238 398
use T_flip_flop  T_flip_flop_0 ~/Desktop/Fossi_cochlea/cochlea_sky130/mag/T_flip_flop
timestamp 1639940534
transform 1 0 -786 0 1 716
box 786 -716 3080 714
use sky130_fd_sc_lp__and2_1  sky130_fd_sc_lp__and2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform -1 0 624 0 -1 715
box -38 -49 518 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 1584 0 -1 715
box -38 -49 710 715
<< end >>
