magic
tech sky130A
magscale 1 2
timestamp 1640489172
<< nwell >>
rect 3389 464 3423 498
rect 5485 314 5549 448
<< pwell >>
rect 3919 99 4039 260
<< poly >>
rect 3918 221 3960 259
rect 3918 138 3999 221
rect 3918 125 3960 138
<< locali >>
rect 3923 221 3964 365
rect 3923 138 3947 221
rect 3999 141 4009 175
rect 3923 102 3964 138
<< viali >>
rect 3389 464 3423 498
rect 3389 382 3423 416
rect 2207 281 2241 315
rect 1872 230 1908 275
rect 3947 138 3999 221
rect 4309 219 4343 253
rect 5670 209 5704 243
rect 5843 206 5878 240
<< metal1 >>
rect 1606 1180 2049 1250
rect 1659 691 1746 730
rect 1971 703 2049 1180
rect 1666 690 1746 691
rect 1714 479 1746 690
rect 3432 650 4045 711
rect 3432 614 4499 650
rect 3886 553 4499 614
rect 5552 551 5644 649
rect 3370 500 3496 523
rect 3370 498 4372 500
rect 1714 435 2238 479
rect 2173 349 2238 435
rect 3370 464 3389 498
rect 3423 464 4372 498
rect 3370 416 4372 464
rect 3370 382 3389 416
rect 3423 382 4372 416
rect 3370 374 4372 382
rect 3370 361 3944 374
rect 4040 361 4372 374
rect 5485 401 5549 448
rect 40 290 1512 330
rect 1467 268 1512 290
rect 1766 275 1931 316
rect 1766 268 1872 275
rect 1467 230 1872 268
rect 1908 230 1931 275
rect 2161 315 2259 349
rect 2161 281 2207 315
rect 2241 281 2259 315
rect 2161 243 2259 281
rect 1467 227 1931 230
rect 1766 192 1931 227
rect 3919 221 4039 260
rect 3919 220 3947 221
rect 3919 138 3946 220
rect 3999 138 4039 221
rect 4255 258 4371 361
rect 5485 343 5926 401
rect 5485 314 5549 343
rect 5601 258 5738 264
rect 4255 253 5738 258
rect 4255 219 4309 253
rect 4343 243 5738 253
rect 4343 219 5670 243
rect 4255 209 5670 219
rect 5704 209 5738 243
rect 4255 205 5738 209
rect 4255 173 4371 205
rect 5601 191 5738 205
rect 5804 240 5926 343
rect 5804 206 5843 240
rect 5878 206 5926 240
rect 5804 189 5926 206
rect 3919 99 4039 138
rect 1650 32 1792 70
rect 1650 -39 1845 32
rect 3457 -17 3762 45
rect 1650 -53 1831 -39
rect 3457 -53 3990 -17
rect 1650 -55 1792 -53
rect 3587 -115 3990 -53
rect 5551 -115 5643 -17
<< via1 >>
rect 87 1019 141 1072
rect 3946 138 3947 220
rect 3947 138 3999 221
<< metal2 >>
rect 62 1086 170 1090
rect 62 1072 4034 1086
rect 62 1019 87 1072
rect 141 1019 4034 1072
rect 62 1016 4034 1019
rect 62 1004 170 1016
rect 3919 221 4034 1016
rect 3919 220 3947 221
rect 3919 138 3946 220
rect 3999 138 4034 221
rect 3919 98 4034 138
use doubletaillatchcomparator  doubletaillatchcomparator_0
timestamp 1640473169
transform 1 0 530 0 1 220
box -540 -220 1140 1030
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640415294
transform 1 0 1826 0 1 -4
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_1
timestamp 1640415294
transform 1 0 3928 0 1 -66
box -38 -49 1670 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 5629 0 1 -66
box -38 -49 710 715
<< end >>
