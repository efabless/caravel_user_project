magic
tech sky130A
magscale 1 2
timestamp 1639959382
<< nwell >>
rect 560 -9313 1121 -8940
<< nsubdiff >>
rect 596 -9204 696 -9182
rect 596 -9238 628 -9204
rect 662 -9238 696 -9204
rect 596 -9260 696 -9238
<< nsubdiffcont >>
rect 628 -9238 662 -9204
<< locali >>
rect 596 -9204 696 -9180
rect 596 -9238 628 -9204
rect 662 -9238 696 -9204
rect 596 -9258 696 -9238
rect 596 -9292 784 -9258
<< metal1 >>
rect 16 1430 60 1432
rect 4 1331 103 1430
rect 2220 1428 2352 1430
rect 2252 1422 2352 1428
rect 2252 1340 2262 1422
rect 2342 1340 2352 1422
rect 2252 1331 2352 1340
rect -82 1286 -14 1292
rect -82 1234 -76 1286
rect -20 1278 -14 1286
rect -20 1244 38 1278
rect -20 1234 -14 1244
rect -82 1228 -14 1234
rect -174 926 -106 932
rect -174 874 -168 926
rect -112 924 -106 926
rect -112 876 4 924
rect -112 874 -106 876
rect -174 868 -106 874
rect 2162 754 2481 764
rect 2162 672 2390 754
rect 2470 672 2481 754
rect 2162 665 2481 672
rect 2260 294 2262 340
rect 2252 88 2352 98
rect 2252 6 2264 88
rect 2344 6 2352 88
rect 2252 -1 2352 6
rect -84 -46 -16 -40
rect -84 -98 -78 -46
rect -22 -54 -16 -46
rect -22 -88 38 -54
rect -22 -98 -16 -88
rect -84 -104 -16 -98
rect -174 -406 -106 -400
rect -174 -458 -168 -406
rect -112 -408 -106 -406
rect -112 -456 4 -408
rect -112 -458 -106 -456
rect -174 -464 -106 -458
rect 2162 -578 2479 -568
rect 2162 -660 2388 -578
rect 2468 -660 2479 -578
rect 2162 -667 2479 -660
rect 2260 -1038 2264 -992
rect 2252 -1244 2352 -1234
rect 2252 -1326 2262 -1244
rect 2342 -1326 2352 -1244
rect 2252 -1333 2352 -1326
rect -84 -1376 -16 -1370
rect -84 -1428 -78 -1376
rect -22 -1386 -16 -1376
rect -22 -1420 38 -1386
rect -22 -1428 -16 -1420
rect -84 -1434 -16 -1428
rect -174 -1738 -106 -1732
rect -174 -1790 -168 -1738
rect -112 -1740 -106 -1738
rect -112 -1788 4 -1740
rect -112 -1790 -106 -1788
rect -174 -1796 -106 -1790
rect 2162 -1908 2479 -1900
rect 2162 -1990 2390 -1908
rect 2470 -1990 2479 -1908
rect 2162 -1999 2479 -1990
rect 2260 -2370 2264 -2324
rect 2252 -2574 2352 -2566
rect 2252 -2656 2264 -2574
rect 2344 -2656 2352 -2574
rect 2252 -2665 2352 -2656
rect -84 -2710 -16 -2704
rect -84 -2762 -78 -2710
rect -22 -2718 -16 -2710
rect -22 -2752 38 -2718
rect -22 -2762 -16 -2752
rect -84 -2768 -16 -2762
rect -174 -3070 -106 -3064
rect -174 -3122 -168 -3070
rect -112 -3072 -106 -3070
rect -112 -3120 4 -3072
rect -112 -3122 -106 -3120
rect -174 -3128 -106 -3122
rect 2162 -3244 2479 -3232
rect 2162 -3326 2388 -3244
rect 2468 -3326 2479 -3244
rect 2162 -3331 2479 -3326
rect 2260 -3702 2264 -3656
rect 2252 -3910 2352 -3898
rect 2252 -3992 2262 -3910
rect 2342 -3992 2352 -3910
rect 2252 -3997 2352 -3992
rect -84 -4042 -16 -4036
rect -84 -4094 -78 -4042
rect -22 -4050 -16 -4042
rect -22 -4084 38 -4050
rect -22 -4094 -16 -4084
rect -84 -4100 -16 -4094
rect -174 -4402 -106 -4396
rect -174 -4454 -168 -4402
rect -112 -4404 -106 -4402
rect -112 -4452 4 -4404
rect -112 -4454 -106 -4452
rect -174 -4460 -106 -4454
rect 2162 -4576 2479 -4564
rect 2162 -4658 2390 -4576
rect 2470 -4658 2479 -4576
rect 2162 -4663 2479 -4658
rect 2260 -5034 2264 -4988
rect 2252 -5238 2352 -5230
rect 2252 -5320 2262 -5238
rect 2342 -5320 2352 -5238
rect 2252 -5329 2352 -5320
rect -84 -5374 -16 -5368
rect -84 -5426 -78 -5374
rect -22 -5382 -16 -5374
rect -22 -5416 38 -5382
rect -22 -5426 -16 -5416
rect -84 -5432 -16 -5426
rect -174 -5734 -106 -5728
rect -174 -5786 -168 -5734
rect -112 -5736 -106 -5734
rect -112 -5784 4 -5736
rect -112 -5786 -106 -5784
rect -174 -5792 -106 -5786
rect 2162 -5904 2479 -5896
rect 2162 -5986 2388 -5904
rect 2468 -5986 2479 -5904
rect 2162 -5995 2479 -5986
rect 2260 -6366 2264 -6320
rect 2252 -6570 2352 -6562
rect 2252 -6652 2264 -6570
rect 2344 -6652 2352 -6570
rect 2252 -6661 2352 -6652
rect -84 -6704 -16 -6698
rect -84 -6756 -78 -6704
rect -22 -6714 -16 -6704
rect -22 -6748 38 -6714
rect -22 -6756 -16 -6748
rect -84 -6762 -16 -6756
rect -174 -7066 -106 -7060
rect -174 -7118 -168 -7066
rect -112 -7068 -106 -7066
rect -112 -7116 4 -7068
rect -112 -7118 -106 -7116
rect -174 -7124 -106 -7118
rect 2162 -7234 2481 -7228
rect 2162 -7316 2390 -7234
rect 2470 -7316 2481 -7234
rect 2162 -7327 2481 -7316
rect 2260 -7698 2266 -7652
rect 2252 -7902 2352 -7894
rect 2252 -7984 2264 -7902
rect 2344 -7984 2352 -7902
rect 2252 -7993 2352 -7984
rect -84 -8038 -16 -8032
rect -84 -8090 -78 -8038
rect -22 -8046 -16 -8038
rect -22 -8080 38 -8046
rect -22 -8090 -16 -8080
rect -84 -8096 -16 -8090
rect 2264 -8360 2270 -8300
rect -174 -8398 -106 -8392
rect -174 -8450 -168 -8398
rect -112 -8400 -106 -8398
rect -112 -8448 38 -8400
rect -112 -8450 -106 -8448
rect -174 -8456 -106 -8450
rect 2162 -8567 2481 -8560
rect 2162 -8649 2392 -8567
rect 2472 -8649 2481 -8567
rect 2162 -8659 2481 -8649
rect 2 -8870 72 -8864
rect 2 -8926 10 -8870
rect 66 -8926 72 -8870
rect 2 -8930 72 -8926
rect 1427 -9235 2352 -9226
rect 1427 -9317 2262 -9235
rect 2342 -9317 2352 -9235
rect 1427 -9324 2352 -9317
<< via1 >>
rect 2262 1340 2342 1422
rect -76 1234 -20 1286
rect -168 874 -112 926
rect 2390 672 2470 754
rect 2264 6 2344 88
rect -78 -98 -22 -46
rect -168 -458 -112 -406
rect 2388 -660 2468 -578
rect 2262 -1326 2342 -1244
rect -78 -1428 -22 -1376
rect -168 -1790 -112 -1738
rect 2390 -1990 2470 -1908
rect 2264 -2656 2344 -2574
rect -78 -2762 -22 -2710
rect -168 -3122 -112 -3070
rect 2388 -3326 2468 -3244
rect 2262 -3992 2342 -3910
rect -78 -4094 -22 -4042
rect -168 -4454 -112 -4402
rect 2390 -4658 2470 -4576
rect 2262 -5320 2342 -5238
rect -78 -5426 -22 -5374
rect -168 -5786 -112 -5734
rect 2388 -5986 2468 -5904
rect 2264 -6652 2344 -6570
rect -78 -6756 -22 -6704
rect -168 -7118 -112 -7066
rect 2390 -7316 2470 -7234
rect 2264 -7984 2344 -7902
rect -78 -8090 -22 -8038
rect -168 -8450 -112 -8398
rect 2392 -8649 2472 -8567
rect 10 -8926 66 -8870
rect 2262 -9317 2342 -9235
<< metal2 >>
rect 16 1430 60 1432
rect -162 932 -118 1430
rect -72 1292 -28 1430
rect 2252 1422 2352 1430
rect 2252 1340 2262 1422
rect 2342 1340 2352 1422
rect -82 1286 -14 1292
rect -82 1234 -76 1286
rect -20 1234 -14 1286
rect -82 1228 -14 1234
rect -174 926 -106 932
rect -174 874 -168 926
rect -112 874 -106 926
rect -174 868 -106 874
rect -162 -400 -118 868
rect -72 -40 -28 1228
rect 2252 88 2352 1340
rect 2252 6 2264 88
rect 2344 6 2352 88
rect -84 -46 -16 -40
rect -84 -98 -78 -46
rect -22 -98 -16 -46
rect -84 -104 -16 -98
rect -174 -406 -106 -400
rect -174 -458 -168 -406
rect -112 -458 -106 -406
rect -174 -464 -106 -458
rect -162 -1732 -118 -464
rect -72 -1370 -28 -104
rect 2252 -1244 2352 6
rect 2252 -1326 2262 -1244
rect 2342 -1326 2352 -1244
rect -84 -1376 -16 -1370
rect -84 -1428 -78 -1376
rect -22 -1428 -16 -1376
rect -84 -1434 -16 -1428
rect -174 -1738 -106 -1732
rect -174 -1790 -168 -1738
rect -112 -1790 -106 -1738
rect -174 -1796 -106 -1790
rect -162 -3064 -118 -1796
rect -72 -2704 -28 -1434
rect 2252 -2574 2352 -1326
rect 2252 -2656 2264 -2574
rect 2344 -2656 2352 -2574
rect -84 -2710 -16 -2704
rect -84 -2762 -78 -2710
rect -22 -2762 -16 -2710
rect -84 -2768 -16 -2762
rect -174 -3070 -106 -3064
rect -174 -3122 -168 -3070
rect -112 -3122 -106 -3070
rect -174 -3128 -106 -3122
rect -162 -4396 -118 -3128
rect -72 -4036 -28 -2768
rect 2252 -3910 2352 -2656
rect 2252 -3992 2262 -3910
rect 2342 -3992 2352 -3910
rect -84 -4042 -16 -4036
rect -84 -4094 -78 -4042
rect -22 -4094 -16 -4042
rect -84 -4100 -16 -4094
rect -174 -4402 -106 -4396
rect -174 -4454 -168 -4402
rect -112 -4454 -106 -4402
rect -174 -4460 -106 -4454
rect -162 -5728 -118 -4460
rect -72 -5368 -28 -4100
rect 2252 -5238 2352 -3992
rect 2252 -5320 2262 -5238
rect 2342 -5320 2352 -5238
rect -84 -5374 -16 -5368
rect -84 -5426 -78 -5374
rect -22 -5426 -16 -5374
rect -84 -5432 -16 -5426
rect -174 -5734 -106 -5728
rect -174 -5786 -168 -5734
rect -112 -5786 -106 -5734
rect -174 -5792 -106 -5786
rect -162 -7060 -118 -5792
rect -72 -6698 -28 -5432
rect 2252 -6570 2352 -5320
rect 2252 -6652 2264 -6570
rect 2344 -6652 2352 -6570
rect -84 -6704 -16 -6698
rect -84 -6756 -78 -6704
rect -22 -6756 -16 -6704
rect -84 -6762 -16 -6756
rect -174 -7066 -106 -7060
rect -174 -7118 -168 -7066
rect -112 -7118 -106 -7066
rect -174 -7124 -106 -7118
rect -162 -8392 -118 -7124
rect -72 -8032 -28 -6762
rect -84 -8038 -16 -8032
rect -84 -8090 -78 -8038
rect -22 -8090 -16 -8038
rect -84 -8096 -16 -8090
rect -174 -8398 -106 -8392
rect -174 -8450 -168 -8398
rect -112 -8450 -106 -8398
rect -174 -8456 -106 -8450
rect 16 -8864 60 -7844
rect 2150 -8344 2202 -7830
rect 2252 -7902 2352 -6652
rect 2252 -7984 2264 -7902
rect 2344 -7984 2352 -7902
rect 2 -8870 72 -8864
rect 2 -8926 10 -8870
rect 66 -8926 72 -8870
rect 2 -8930 72 -8926
rect 2252 -9235 2352 -7984
rect 2382 754 2480 1430
rect 2382 672 2390 754
rect 2470 672 2480 754
rect 2382 -578 2480 672
rect 2382 -660 2388 -578
rect 2468 -660 2480 -578
rect 2382 -1908 2480 -660
rect 2382 -1990 2390 -1908
rect 2470 -1990 2480 -1908
rect 2382 -3244 2480 -1990
rect 2382 -3326 2388 -3244
rect 2468 -3326 2480 -3244
rect 2382 -4576 2480 -3326
rect 2382 -4658 2390 -4576
rect 2470 -4658 2480 -4576
rect 2382 -5904 2480 -4658
rect 2382 -5986 2388 -5904
rect 2468 -5986 2480 -5904
rect 2382 -7234 2480 -5986
rect 2382 -7316 2390 -7234
rect 2470 -7316 2480 -7234
rect 2382 -8567 2480 -7316
rect 2382 -8649 2392 -8567
rect 2472 -8649 2480 -8567
rect 2382 -8659 2480 -8649
rect 2252 -9317 2262 -9235
rect 2342 -9317 2352 -9235
rect 2252 -9322 2352 -9317
use asyn_gr_counter_cell  asyn_gr_counter_cell_2
timestamp 1639940697
transform 1 0 2 0 1 -2664
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_1
timestamp 1639940697
transform 1 0 2 0 1 -1332
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_0
timestamp 1639940697
transform 1 0 2 0 1 0
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_6
timestamp 1639940697
transform 1 0 2 0 1 -7992
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_5
timestamp 1639940697
transform 1 0 2 0 1 -6660
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_4
timestamp 1639940697
transform 1 0 2 0 1 -5328
box -32 0 2262 1430
use asyn_gr_counter_cell  asyn_gr_counter_cell_3
timestamp 1639940697
transform 1 0 2 0 1 -3996
box -32 0 2262 1430
use T_flip_flop  T_flip_flop_0
timestamp 1639940534
transform 1 0 -816 0 1 -8608
box 786 -716 3080 714
<< labels >>
rlabel metal2 -52 1430 -52 1430 1 RSTB
port 1 n
rlabel metal2 -144 1430 -144 1430 1 CLK
port 3 n
rlabel metal1 2260 314 2260 314 3 Q0
port 4 e
rlabel metal1 2260 -1016 2260 -1016 3 Q1
port 5 e
rlabel metal1 2260 -2352 2260 -2352 3 Q2
port 6 e
rlabel metal1 2260 -3680 2260 -3680 3 Q3
port 7 e
rlabel metal1 2260 -5016 2260 -5016 3 Q4
port 8 e
rlabel metal1 2260 -6346 2260 -6346 3 Q5
port 9 e
rlabel metal1 2260 -7678 2260 -7678 3 Q6
port 10 e
rlabel metal1 2264 -8334 2264 -8334 3 Q7
port 11 e
rlabel metal2 36 1432 36 1432 1 EN
port 2 n
rlabel metal2 2300 1430 2300 1430 1 Vdd
port 12 n
rlabel metal2 2430 1430 2430 1430 1 gnd
port 13 n
<< end >>
