magic
tech sky130A
magscale 1 2
timestamp 1640506818
<< nwell >>
rect 1058 702 1722 998
<< poly >>
rect 1178 1028 1208 1098
<< locali >>
rect 3242 618 3282 664
<< viali >>
rect 4874 626 4914 670
rect 1718 432 1758 478
rect 2030 470 2076 524
rect 3344 440 3380 480
rect 3656 468 3700 522
rect 4994 468 5034 526
rect 5162 442 5196 476
rect 3244 326 3282 372
<< metal1 >>
rect 1536 1162 2002 1232
rect 28 862 68 1010
rect 1916 914 2002 1162
rect 28 822 1598 862
rect 1558 724 1598 822
rect 1558 684 3410 724
rect 1584 558 2094 592
rect 1584 552 2096 558
rect 2004 524 2096 552
rect 1696 478 1768 524
rect 1414 438 1718 478
rect 1414 312 1452 438
rect 1696 432 1718 438
rect 1758 432 1768 478
rect 2004 470 2030 524
rect 2076 470 2096 524
rect 2004 442 2096 470
rect 3332 480 3410 684
rect 4860 670 4930 746
rect 4860 626 4874 670
rect 4914 626 4930 670
rect 4860 582 4930 626
rect 3332 440 3344 480
rect 3380 440 3410 480
rect 1696 368 1768 432
rect 3232 372 3292 434
rect 3332 382 3410 440
rect 3628 522 3730 558
rect 3628 468 3656 522
rect 3700 468 3730 522
rect 452 272 1452 312
rect 3232 326 3244 372
rect 3282 342 3292 372
rect 3628 342 3730 468
rect 4860 526 5042 582
rect 4860 468 4994 526
rect 5034 468 5042 526
rect 4860 446 5042 468
rect 5134 476 5216 490
rect 5134 442 5162 476
rect 5196 442 5216 476
rect 5134 342 5216 442
rect 3282 326 5216 342
rect 3232 280 5216 326
rect 1934 52 2020 166
rect 1598 -18 2020 52
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 4944 0 1 200
box -38 -49 710 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_1 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640415294
transform 1 0 3312 0 1 200
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_0
timestamp 1640415294
transform 1 0 1680 0 1 200
box -38 -49 1670 715
use doubletaillatchcomparator  doubletaillatchcomparator_0 ~/fossi_cochlea/mag/comparator
timestamp 1640503333
transform 1 0 488 0 1 202
box -540 -220 1140 1030
<< end >>
