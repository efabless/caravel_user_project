magic
tech sky130A
magscale 1 2
timestamp 1621087811
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 106 960 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10138 119200 10194 120000
rect 11702 119200 11758 120000
rect 13266 119200 13322 120000
rect 14830 119200 14886 120000
rect 16394 119200 16450 120000
rect 17958 119200 18014 120000
rect 19522 119200 19578 120000
rect 21086 119200 21142 120000
rect 22650 119200 22706 120000
rect 24214 119200 24270 120000
rect 25778 119200 25834 120000
rect 27342 119200 27398 120000
rect 28906 119200 28962 120000
rect 30470 119200 30526 120000
rect 32034 119200 32090 120000
rect 33598 119200 33654 120000
rect 35162 119200 35218 120000
rect 36726 119200 36782 120000
rect 38290 119200 38346 120000
rect 39854 119200 39910 120000
rect 41418 119200 41474 120000
rect 42982 119200 43038 120000
rect 44546 119200 44602 120000
rect 46110 119200 46166 120000
rect 47674 119200 47730 120000
rect 49238 119200 49294 120000
rect 50802 119200 50858 120000
rect 52366 119200 52422 120000
rect 53930 119200 53986 120000
rect 55494 119200 55550 120000
rect 57058 119200 57114 120000
rect 58622 119200 58678 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63314 119200 63370 120000
rect 64878 119200 64934 120000
rect 66442 119200 66498 120000
rect 68006 119200 68062 120000
rect 69570 119200 69626 120000
rect 71134 119200 71190 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75826 119200 75882 120000
rect 77390 119200 77446 120000
rect 78954 119200 79010 120000
rect 80518 119200 80574 120000
rect 82082 119200 82138 120000
rect 83646 119200 83702 120000
rect 85210 119200 85266 120000
rect 86774 119200 86830 120000
rect 88338 119200 88394 120000
rect 89902 119200 89958 120000
rect 91558 119200 91614 120000
rect 93122 119200 93178 120000
rect 94686 119200 94742 120000
rect 96250 119200 96306 120000
rect 97814 119200 97870 120000
rect 99378 119200 99434 120000
rect 100942 119200 100998 120000
rect 102506 119200 102562 120000
rect 104070 119200 104126 120000
rect 105634 119200 105690 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110326 119200 110382 120000
rect 111890 119200 111946 120000
rect 113454 119200 113510 120000
rect 115018 119200 115074 120000
rect 116582 119200 116638 120000
rect 118146 119200 118202 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122838 119200 122894 120000
rect 124402 119200 124458 120000
rect 125966 119200 126022 120000
rect 127530 119200 127586 120000
rect 129094 119200 129150 120000
rect 130658 119200 130714 120000
rect 132222 119200 132278 120000
rect 133786 119200 133842 120000
rect 135350 119200 135406 120000
rect 136914 119200 136970 120000
rect 138478 119200 138534 120000
rect 140042 119200 140098 120000
rect 141606 119200 141662 120000
rect 143170 119200 143226 120000
rect 144734 119200 144790 120000
rect 146298 119200 146354 120000
rect 147862 119200 147918 120000
rect 149426 119200 149482 120000
rect 150990 119200 151046 120000
rect 152554 119200 152610 120000
rect 154118 119200 154174 120000
rect 155682 119200 155738 120000
rect 157246 119200 157302 120000
rect 158810 119200 158866 120000
rect 160374 119200 160430 120000
rect 161938 119200 161994 120000
rect 163502 119200 163558 120000
rect 165066 119200 165122 120000
rect 166630 119200 166686 120000
rect 168194 119200 168250 120000
rect 169758 119200 169814 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119200
rect 866 119144 2262 119200
rect 2430 119144 3826 119200
rect 3994 119144 5390 119200
rect 5558 119144 6954 119200
rect 7122 119144 8518 119200
rect 8686 119144 10082 119200
rect 10250 119144 11646 119200
rect 11814 119144 13210 119200
rect 13378 119144 14774 119200
rect 14942 119144 16338 119200
rect 16506 119144 17902 119200
rect 18070 119144 19466 119200
rect 19634 119144 21030 119200
rect 21198 119144 22594 119200
rect 22762 119144 24158 119200
rect 24326 119144 25722 119200
rect 25890 119144 27286 119200
rect 27454 119144 28850 119200
rect 29018 119144 30414 119200
rect 30582 119144 31978 119200
rect 32146 119144 33542 119200
rect 33710 119144 35106 119200
rect 35274 119144 36670 119200
rect 36838 119144 38234 119200
rect 38402 119144 39798 119200
rect 39966 119144 41362 119200
rect 41530 119144 42926 119200
rect 43094 119144 44490 119200
rect 44658 119144 46054 119200
rect 46222 119144 47618 119200
rect 47786 119144 49182 119200
rect 49350 119144 50746 119200
rect 50914 119144 52310 119200
rect 52478 119144 53874 119200
rect 54042 119144 55438 119200
rect 55606 119144 57002 119200
rect 57170 119144 58566 119200
rect 58734 119144 60130 119200
rect 60298 119144 61694 119200
rect 61862 119144 63258 119200
rect 63426 119144 64822 119200
rect 64990 119144 66386 119200
rect 66554 119144 67950 119200
rect 68118 119144 69514 119200
rect 69682 119144 71078 119200
rect 71246 119144 72642 119200
rect 72810 119144 74206 119200
rect 74374 119144 75770 119200
rect 75938 119144 77334 119200
rect 77502 119144 78898 119200
rect 79066 119144 80462 119200
rect 80630 119144 82026 119200
rect 82194 119144 83590 119200
rect 83758 119144 85154 119200
rect 85322 119144 86718 119200
rect 86886 119144 88282 119200
rect 88450 119144 89846 119200
rect 90014 119144 91502 119200
rect 91670 119144 93066 119200
rect 93234 119144 94630 119200
rect 94798 119144 96194 119200
rect 96362 119144 97758 119200
rect 97926 119144 99322 119200
rect 99490 119144 100886 119200
rect 101054 119144 102450 119200
rect 102618 119144 104014 119200
rect 104182 119144 105578 119200
rect 105746 119144 107142 119200
rect 107310 119144 108706 119200
rect 108874 119144 110270 119200
rect 110438 119144 111834 119200
rect 112002 119144 113398 119200
rect 113566 119144 114962 119200
rect 115130 119144 116526 119200
rect 116694 119144 118090 119200
rect 118258 119144 119654 119200
rect 119822 119144 121218 119200
rect 121386 119144 122782 119200
rect 122950 119144 124346 119200
rect 124514 119144 125910 119200
rect 126078 119144 127474 119200
rect 127642 119144 129038 119200
rect 129206 119144 130602 119200
rect 130770 119144 132166 119200
rect 132334 119144 133730 119200
rect 133898 119144 135294 119200
rect 135462 119144 136858 119200
rect 137026 119144 138422 119200
rect 138590 119144 139986 119200
rect 140154 119144 141550 119200
rect 141718 119144 143114 119200
rect 143282 119144 144678 119200
rect 144846 119144 146242 119200
rect 146410 119144 147806 119200
rect 147974 119144 149370 119200
rect 149538 119144 150934 119200
rect 151102 119144 152498 119200
rect 152666 119144 154062 119200
rect 154230 119144 155626 119200
rect 155794 119144 157190 119200
rect 157358 119144 158754 119200
rect 158922 119144 160318 119200
rect 160486 119144 161882 119200
rect 162050 119144 163446 119200
rect 163614 119144 165010 119200
rect 165178 119144 166574 119200
rect 166742 119144 168138 119200
rect 168306 119144 169702 119200
rect 169870 119144 171266 119200
rect 171434 119144 172830 119200
rect 172998 119144 174394 119200
rect 174562 119144 175958 119200
rect 176126 119144 177522 119200
rect 177690 119144 179086 119200
rect 179254 119144 179840 119200
rect 112 856 179840 119144
rect 222 800 330 856
rect 498 800 698 856
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4378 856
rect 4546 800 4746 856
rect 4914 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5850 856
rect 6018 800 6218 856
rect 6386 800 6586 856
rect 6754 800 6954 856
rect 7122 800 7322 856
rect 7490 800 7690 856
rect 7858 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8794 856
rect 8962 800 9162 856
rect 9330 800 9530 856
rect 9698 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10634 856
rect 10802 800 11002 856
rect 11170 800 11370 856
rect 11538 800 11738 856
rect 11906 800 12106 856
rect 12274 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13578 856
rect 13746 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15050 856
rect 15218 800 15418 856
rect 15586 800 15786 856
rect 15954 800 16154 856
rect 16322 800 16522 856
rect 16690 800 16890 856
rect 17058 800 17258 856
rect 17426 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18730 856
rect 18898 800 19098 856
rect 19266 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23146 856
rect 23314 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 26090 856
rect 26258 800 26458 856
rect 26626 800 26826 856
rect 26994 800 27194 856
rect 27362 800 27562 856
rect 27730 800 27930 856
rect 28098 800 28298 856
rect 28466 800 28666 856
rect 28834 800 29034 856
rect 29202 800 29402 856
rect 29570 800 29770 856
rect 29938 800 30138 856
rect 30306 800 30506 856
rect 30674 800 30874 856
rect 31042 800 31242 856
rect 31410 800 31610 856
rect 31778 800 31978 856
rect 32146 800 32346 856
rect 32514 800 32714 856
rect 32882 800 33082 856
rect 33250 800 33450 856
rect 33618 800 33818 856
rect 33986 800 34186 856
rect 34354 800 34554 856
rect 34722 800 34922 856
rect 35090 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38234 856
rect 38402 800 38602 856
rect 38770 800 38970 856
rect 39138 800 39338 856
rect 39506 800 39706 856
rect 39874 800 40074 856
rect 40242 800 40442 856
rect 40610 800 40810 856
rect 40978 800 41178 856
rect 41346 800 41546 856
rect 41714 800 41914 856
rect 42082 800 42282 856
rect 42450 800 42650 856
rect 42818 800 43018 856
rect 43186 800 43386 856
rect 43554 800 43754 856
rect 43922 800 44122 856
rect 44290 800 44490 856
rect 44658 800 44858 856
rect 45026 800 45226 856
rect 45394 800 45594 856
rect 45762 800 45962 856
rect 46130 800 46330 856
rect 46498 800 46698 856
rect 46866 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47802 856
rect 47970 800 48170 856
rect 48338 800 48538 856
rect 48706 800 48906 856
rect 49074 800 49274 856
rect 49442 800 49642 856
rect 49810 800 50010 856
rect 50178 800 50378 856
rect 50546 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51482 856
rect 51650 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52586 856
rect 52754 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53690 856
rect 53858 800 54058 856
rect 54226 800 54426 856
rect 54594 800 54794 856
rect 54962 800 55162 856
rect 55330 800 55530 856
rect 55698 800 55898 856
rect 56066 800 56266 856
rect 56434 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57738 856
rect 57906 800 58106 856
rect 58274 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59210 856
rect 59378 800 59578 856
rect 59746 800 59946 856
rect 60114 800 60222 856
rect 60390 800 60590 856
rect 60758 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61694 856
rect 61862 800 62062 856
rect 62230 800 62430 856
rect 62598 800 62798 856
rect 62966 800 63166 856
rect 63334 800 63534 856
rect 63702 800 63902 856
rect 64070 800 64270 856
rect 64438 800 64638 856
rect 64806 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65742 856
rect 65910 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66846 856
rect 67014 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68318 856
rect 68486 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69422 856
rect 69590 800 69790 856
rect 69958 800 70158 856
rect 70326 800 70526 856
rect 70694 800 70894 856
rect 71062 800 71262 856
rect 71430 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73838 856
rect 74006 800 74206 856
rect 74374 800 74574 856
rect 74742 800 74942 856
rect 75110 800 75310 856
rect 75478 800 75678 856
rect 75846 800 76046 856
rect 76214 800 76414 856
rect 76582 800 76782 856
rect 76950 800 77150 856
rect 77318 800 77518 856
rect 77686 800 77886 856
rect 78054 800 78254 856
rect 78422 800 78622 856
rect 78790 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79726 856
rect 79894 800 80094 856
rect 80262 800 80462 856
rect 80630 800 80830 856
rect 80998 800 81198 856
rect 81366 800 81566 856
rect 81734 800 81934 856
rect 82102 800 82302 856
rect 82470 800 82670 856
rect 82838 800 83038 856
rect 83206 800 83406 856
rect 83574 800 83774 856
rect 83942 800 84142 856
rect 84310 800 84510 856
rect 84678 800 84878 856
rect 85046 800 85246 856
rect 85414 800 85614 856
rect 85782 800 85982 856
rect 86150 800 86350 856
rect 86518 800 86718 856
rect 86886 800 87086 856
rect 87254 800 87454 856
rect 87622 800 87822 856
rect 87990 800 88190 856
rect 88358 800 88558 856
rect 88726 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90398 856
rect 90566 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92606 856
rect 92774 800 92974 856
rect 93142 800 93342 856
rect 93510 800 93710 856
rect 93878 800 94078 856
rect 94246 800 94446 856
rect 94614 800 94814 856
rect 94982 800 95182 856
rect 95350 800 95550 856
rect 95718 800 95918 856
rect 96086 800 96286 856
rect 96454 800 96654 856
rect 96822 800 97022 856
rect 97190 800 97390 856
rect 97558 800 97758 856
rect 97926 800 98126 856
rect 98294 800 98494 856
rect 98662 800 98862 856
rect 99030 800 99230 856
rect 99398 800 99598 856
rect 99766 800 99966 856
rect 100134 800 100334 856
rect 100502 800 100702 856
rect 100870 800 101070 856
rect 101238 800 101438 856
rect 101606 800 101806 856
rect 101974 800 102174 856
rect 102342 800 102542 856
rect 102710 800 102910 856
rect 103078 800 103278 856
rect 103446 800 103646 856
rect 103814 800 104014 856
rect 104182 800 104382 856
rect 104550 800 104750 856
rect 104918 800 105118 856
rect 105286 800 105486 856
rect 105654 800 105854 856
rect 106022 800 106222 856
rect 106390 800 106590 856
rect 106758 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107694 856
rect 107862 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108798 856
rect 108966 800 109166 856
rect 109334 800 109534 856
rect 109702 800 109902 856
rect 110070 800 110270 856
rect 110438 800 110638 856
rect 110806 800 111006 856
rect 111174 800 111374 856
rect 111542 800 111742 856
rect 111910 800 112110 856
rect 112278 800 112478 856
rect 112646 800 112846 856
rect 113014 800 113214 856
rect 113382 800 113582 856
rect 113750 800 113950 856
rect 114118 800 114318 856
rect 114486 800 114686 856
rect 114854 800 115054 856
rect 115222 800 115422 856
rect 115590 800 115790 856
rect 115958 800 116158 856
rect 116326 800 116526 856
rect 116694 800 116894 856
rect 117062 800 117262 856
rect 117430 800 117630 856
rect 117798 800 117998 856
rect 118166 800 118366 856
rect 118534 800 118734 856
rect 118902 800 119102 856
rect 119270 800 119470 856
rect 119638 800 119838 856
rect 120006 800 120114 856
rect 120282 800 120482 856
rect 120650 800 120850 856
rect 121018 800 121218 856
rect 121386 800 121586 856
rect 121754 800 121954 856
rect 122122 800 122322 856
rect 122490 800 122690 856
rect 122858 800 123058 856
rect 123226 800 123426 856
rect 123594 800 123794 856
rect 123962 800 124162 856
rect 124330 800 124530 856
rect 124698 800 124898 856
rect 125066 800 125266 856
rect 125434 800 125634 856
rect 125802 800 126002 856
rect 126170 800 126370 856
rect 126538 800 126738 856
rect 126906 800 127106 856
rect 127274 800 127474 856
rect 127642 800 127842 856
rect 128010 800 128210 856
rect 128378 800 128578 856
rect 128746 800 128946 856
rect 129114 800 129314 856
rect 129482 800 129682 856
rect 129850 800 130050 856
rect 130218 800 130418 856
rect 130586 800 130786 856
rect 130954 800 131154 856
rect 131322 800 131522 856
rect 131690 800 131890 856
rect 132058 800 132258 856
rect 132426 800 132626 856
rect 132794 800 132994 856
rect 133162 800 133362 856
rect 133530 800 133730 856
rect 133898 800 134098 856
rect 134266 800 134466 856
rect 134634 800 134834 856
rect 135002 800 135202 856
rect 135370 800 135570 856
rect 135738 800 135938 856
rect 136106 800 136306 856
rect 136474 800 136674 856
rect 136842 800 137042 856
rect 137210 800 137410 856
rect 137578 800 137778 856
rect 137946 800 138146 856
rect 138314 800 138514 856
rect 138682 800 138882 856
rect 139050 800 139250 856
rect 139418 800 139618 856
rect 139786 800 139986 856
rect 140154 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141090 856
rect 141258 800 141458 856
rect 141626 800 141826 856
rect 141994 800 142194 856
rect 142362 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143298 856
rect 143466 800 143666 856
rect 143834 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145874 856
rect 146042 800 146242 856
rect 146410 800 146610 856
rect 146778 800 146978 856
rect 147146 800 147346 856
rect 147514 800 147714 856
rect 147882 800 148082 856
rect 148250 800 148450 856
rect 148618 800 148818 856
rect 148986 800 149186 856
rect 149354 800 149554 856
rect 149722 800 149922 856
rect 150090 800 150290 856
rect 150458 800 150658 856
rect 150826 800 151026 856
rect 151194 800 151394 856
rect 151562 800 151762 856
rect 151930 800 152130 856
rect 152298 800 152498 856
rect 152666 800 152866 856
rect 153034 800 153234 856
rect 153402 800 153602 856
rect 153770 800 153970 856
rect 154138 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160594 856
rect 160762 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162066 856
rect 162234 800 162434 856
rect 162602 800 162802 856
rect 162970 800 163170 856
rect 163338 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164274 856
rect 164442 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166482 856
rect 166650 800 166850 856
rect 167018 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167954 856
rect 168122 800 168322 856
rect 168490 800 168690 856
rect 168858 800 169058 856
rect 169226 800 169426 856
rect 169594 800 169794 856
rect 169962 800 170162 856
rect 170330 800 170530 856
rect 170698 800 170898 856
rect 171066 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173106 856
rect 173274 800 173474 856
rect 173642 800 173842 856
rect 174010 800 174210 856
rect 174378 800 174578 856
rect 174746 800 174946 856
rect 175114 800 175314 856
rect 175482 800 175682 856
rect 175850 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178258 856
rect 178426 800 178626 856
rect 178794 800 178994 856
rect 179162 800 179362 856
rect 179530 800 179730 856
<< metal3 >>
rect 0 59984 800 60104
rect 179200 59984 180000 60104
<< obsm3 >>
rect 800 60184 179200 117537
rect 880 59904 179120 60184
rect 800 1939 179200 59904
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 8339 2048 19488 52869
rect 19968 2096 20148 52869
rect 20628 2096 20808 52869
rect 21288 2096 21468 52869
rect 21948 2096 34848 52869
rect 19968 2048 34848 2096
rect 35328 2096 35508 52869
rect 35988 2096 36168 52869
rect 36648 2096 36828 52869
rect 37308 2096 50208 52869
rect 35328 2048 50208 2096
rect 50688 2096 50868 52869
rect 51348 2096 51528 52869
rect 52008 2096 52188 52869
rect 52668 2096 65568 52869
rect 50688 2048 65568 2096
rect 66048 2096 66228 52869
rect 66708 2096 66888 52869
rect 67368 2096 67548 52869
rect 68028 2096 80928 52869
rect 66048 2048 80928 2096
rect 81408 2096 81588 52869
rect 82068 2096 82248 52869
rect 82728 2096 82908 52869
rect 83388 2096 96288 52869
rect 81408 2048 96288 2096
rect 96768 2096 96948 52869
rect 97428 2096 97608 52869
rect 98088 2096 98268 52869
rect 98748 2096 105090 52869
rect 96768 2048 105090 2096
rect 8339 1939 105090 2048
<< obsm5 >>
rect 68012 36220 105132 46740
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52366 119200 52422 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57058 119200 57114 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 66442 119200 66498 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71134 119200 71190 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 75826 119200 75882 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 85210 119200 85266 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 94686 119200 94742 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 99378 119200 99434 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104070 119200 104126 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 113454 119200 113510 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 122838 119200 122894 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 127530 119200 127586 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132222 119200 132278 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10138 119200 10194 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 141606 119200 141662 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 146298 119200 146354 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 150990 119200 151046 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165066 119200 165122 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 174450 119200 174506 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14830 119200 14886 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19522 119200 19578 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 28906 119200 28962 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33598 119200 33654 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38290 119200 38346 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 42982 119200 43038 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49238 119200 49294 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63314 119200 63370 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68006 119200 68062 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 72698 119200 72754 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 77390 119200 77446 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82082 119200 82138 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 86774 119200 86830 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 91558 119200 91614 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 100942 119200 100998 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 110326 119200 110382 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115018 119200 115074 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 124402 119200 124458 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129094 119200 129150 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 133786 119200 133842 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 138478 119200 138534 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11702 119200 11758 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143170 119200 143226 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 147862 119200 147918 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 152554 119200 152610 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157246 119200 157302 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 161938 119200 161994 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 166630 119200 166686 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 171322 119200 171378 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176014 119200 176070 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16394 119200 16450 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21086 119200 21142 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35162 119200 35218 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 39854 119200 39910 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 50802 119200 50858 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 64878 119200 64934 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 78954 119200 79010 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 83646 119200 83702 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 88338 119200 88394 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93122 119200 93178 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 97814 119200 97870 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 102506 119200 102562 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 116582 119200 116638 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 121274 119200 121330 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 125966 119200 126022 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 130658 119200 130714 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 135350 119200 135406 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140042 119200 140098 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13266 119200 13322 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 144734 119200 144790 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 149426 119200 149482 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154118 119200 154174 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 158810 119200 158866 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 163502 119200 163558 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168194 119200 168250 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 172886 119200 172942 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 17958 119200 18014 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22650 119200 22706 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27342 119200 27398 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32034 119200 32090 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 36726 119200 36782 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41418 119200 41474 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46110 119200 46166 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 179142 119200 179198 120000 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179200 59984 180000 60104 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj.gds
string GDS_END 11781276
string GDS_START 498308
<< end >>

