`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***

//***Module***
module register_data #(
        parameter integer WORD_SIZE = 32,
        parameter integer REGISTERS = 32,
        parameter integer LINE_SIZE = 128,
        parameter integer ALUOP_SIZE = 4,
        parameter integer REGDIRSIZE = 5,
        parameter integer ECCBITS = 7
    )
    (
        input  rst_i ,
        input  [WORD_SIZE - 1 : 0] data_to_register_i ,
        input  [REGDIRSIZE - 1 : 0] register_i ,
        input  wregister_i ,
        input  rregister_i ,
        input  [ECCBITS - 1 : 0] parity_bits_i ,
        output reg [WORD_SIZE - 1 : 0] store_data_o ,
        output reg [ECCBITS - 1 : 0] parity_bits_o 
    );

//***Internal logic generated by compiler***  


//***Dumped Internal logic***
    // register bank
    reg [WORD_SIZE + ECCBITS -1:0] r[0:REGISTERS-1];
    wire [ECCBITS - 1:0] parity_bits;

    assign  parity_bits[0] =  parity_bits_i[0];
    assign  parity_bits[1] =  parity_bits_i[1];
    assign  parity_bits[2] =  parity_bits_i[2];
    assign  parity_bits[3] =  parity_bits_i[3];
    assign  parity_bits[4] =  parity_bits_i[4];
    assign  parity_bits[5] =  parity_bits_i[5];
    assign  parity_bits[6] =  parity_bits_i[6] ^ parity_bits_i[0] ^ parity_bits_i[1] ^ parity_bits_i[2] ^ parity_bits_i[3] ^ parity_bits_i[4] ^ parity_bits_i[5]  ; 
    //request
    always @(*) begin
        // calculate last parity bit
        if (rst_i) begin

            r[0] = {WORD_SIZE + ECCBITS{1'b0}};
            r[1] = {WORD_SIZE + ECCBITS{1'b0}};
            r[2] = {WORD_SIZE + ECCBITS{1'b0}};
            r[3] = {WORD_SIZE + ECCBITS{1'b0}};
            r[4] = {WORD_SIZE + ECCBITS{1'b0}};
            r[5] = {WORD_SIZE + ECCBITS{1'b0}};
            r[6] = {WORD_SIZE + ECCBITS{1'b0}};
            r[7] = {WORD_SIZE + ECCBITS{1'b0}};
            /*r[8] = {WORD_SIZE + ECCBITS{1'b0}};
            r[9] = {WORD_SIZE + ECCBITS{1'b0}};
            r[10] = {WORD_SIZE + ECCBITS{1'b0}};
            r[11] = {WORD_SIZE + ECCBITS{1'b0}};
            r[12] = {WORD_SIZE + ECCBITS{1'b0}};
            r[13] = {WORD_SIZE + ECCBITS{1'b0}};
            r[14] = {WORD_SIZE + ECCBITS{1'b0}};
            r[15] = {WORD_SIZE + ECCBITS{1'b0}};*/
           
            store_data_o = {WORD_SIZE}; 
            parity_bits_o = {ECCBITS {1'b0}};
        end
        else if (rregister_i) begin
            store_data_o = r[register_i][WORD_SIZE -1:0];
            parity_bits_o = r[register_i][WORD_SIZE + ECCBITS -1: WORD_SIZE];
        end
        else if (wregister_i) begin
            // calculate parity bits
            r[register_i] = {parity_bits, data_to_register_i};
            store_data_o = {WORD_SIZE {1'b0}}; 
            parity_bits_o = {ECCBITS {1'b0}};
        end 
    end

   
    
//***Handcrafted Internal logic*** 
//TODO
endmodule
