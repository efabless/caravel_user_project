magic
tech sky130A
magscale 1 2
timestamp 1640103014
<< locali >>
rect 67557 57579 67591 57885
rect 72525 56967 72559 57885
rect 106197 57715 106231 57885
rect 301237 57681 301421 57715
rect 301237 57647 301271 57681
rect 383577 57647 383611 57885
rect 238217 57375 238251 57613
rect 344017 57171 344051 57545
rect 364441 57171 364475 57613
rect 384313 57171 384347 57477
rect 449449 57375 449483 57545
rect 464629 57511 464663 57749
rect 446045 57171 446079 57341
rect 468493 57171 468527 57749
rect 275293 56899 275327 57137
rect 471805 57103 471839 57545
rect 390385 6137 390569 6171
rect 390385 6103 390419 6137
rect 347605 5695 347639 6069
rect 389189 5831 389223 6001
rect 392869 5559 392903 6273
rect 393973 5559 394007 6205
rect 282285 5015 282319 5117
rect 272533 4743 272567 4845
rect 282193 4607 282227 4981
rect 282377 4199 282411 5117
rect 134533 3757 134751 3791
rect 134533 3723 134567 3757
rect 134625 3519 134659 3689
rect 134717 3519 134751 3757
rect 135177 3451 135211 3485
rect 135177 3417 135545 3451
rect 151921 2907 151955 3961
rect 451933 3723 451967 3825
rect 451933 3689 452209 3723
rect 454451 3689 455429 3723
rect 461317 3655 461351 3825
rect 498393 3655 498427 3757
rect 160109 3383 160143 3553
rect 430589 3043 430623 3621
rect 461409 3451 461443 3621
<< viali >>
rect 67557 57885 67591 57919
rect 67557 57545 67591 57579
rect 72525 57885 72559 57919
rect 106197 57885 106231 57919
rect 383577 57885 383611 57919
rect 106197 57681 106231 57715
rect 301421 57681 301455 57715
rect 238217 57613 238251 57647
rect 301237 57613 301271 57647
rect 364441 57613 364475 57647
rect 383577 57613 383611 57647
rect 464629 57749 464663 57783
rect 238217 57341 238251 57375
rect 344017 57545 344051 57579
rect 72525 56933 72559 56967
rect 275293 57137 275327 57171
rect 344017 57137 344051 57171
rect 449449 57545 449483 57579
rect 364441 57137 364475 57171
rect 384313 57477 384347 57511
rect 464629 57477 464663 57511
rect 468493 57749 468527 57783
rect 384313 57137 384347 57171
rect 446045 57341 446079 57375
rect 449449 57341 449483 57375
rect 446045 57137 446079 57171
rect 468493 57137 468527 57171
rect 471805 57545 471839 57579
rect 471805 57069 471839 57103
rect 275293 56865 275327 56899
rect 392869 6273 392903 6307
rect 390569 6137 390603 6171
rect 347605 6069 347639 6103
rect 390385 6069 390419 6103
rect 389189 6001 389223 6035
rect 389189 5797 389223 5831
rect 347605 5661 347639 5695
rect 392869 5525 392903 5559
rect 393973 6205 394007 6239
rect 393973 5525 394007 5559
rect 282285 5117 282319 5151
rect 282193 4981 282227 5015
rect 282285 4981 282319 5015
rect 282377 5117 282411 5151
rect 272533 4845 272567 4879
rect 272533 4709 272567 4743
rect 282193 4573 282227 4607
rect 282377 4165 282411 4199
rect 151921 3961 151955 3995
rect 134533 3689 134567 3723
rect 134625 3689 134659 3723
rect 134625 3485 134659 3519
rect 134717 3485 134751 3519
rect 135177 3485 135211 3519
rect 135545 3417 135579 3451
rect 451933 3825 451967 3859
rect 461317 3825 461351 3859
rect 452209 3689 452243 3723
rect 454417 3689 454451 3723
rect 455429 3689 455463 3723
rect 498393 3757 498427 3791
rect 430589 3621 430623 3655
rect 461317 3621 461351 3655
rect 461409 3621 461443 3655
rect 498393 3621 498427 3655
rect 160109 3553 160143 3587
rect 160109 3349 160143 3383
rect 461409 3417 461443 3451
rect 430589 3009 430623 3043
rect 151921 2873 151955 2907
<< metal1 >>
rect 480162 700476 480168 700528
rect 480220 700516 480226 700528
rect 527174 700516 527180 700528
rect 480220 700488 527180 700516
rect 480220 700476 480226 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 402882 700408 402888 700460
rect 402940 700448 402946 700460
rect 429838 700448 429844 700460
rect 402940 700420 429844 700448
rect 402940 700408 402946 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 441522 700408 441528 700460
rect 441580 700448 441586 700460
rect 478506 700448 478512 700460
rect 441580 700420 478512 700448
rect 441580 700408 441586 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 492582 700408 492588 700460
rect 492640 700448 492646 700460
rect 543458 700448 543464 700460
rect 492640 700420 543464 700448
rect 492640 700408 492646 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 378042 700340 378048 700392
rect 378100 700380 378106 700392
rect 397454 700380 397460 700392
rect 378100 700352 397460 700380
rect 378100 700340 378106 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 416682 700340 416688 700392
rect 416740 700380 416746 700392
rect 446122 700380 446128 700392
rect 416740 700352 446128 700380
rect 416740 700340 416746 700352
rect 446122 700340 446128 700352
rect 446180 700340 446186 700392
rect 453942 700340 453948 700392
rect 454000 700380 454006 700392
rect 494790 700380 494796 700392
rect 454000 700352 494796 700380
rect 454000 700340 454006 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 505002 700340 505008 700392
rect 505060 700380 505066 700392
rect 559650 700380 559656 700392
rect 505060 700352 559656 700380
rect 505060 700340 505066 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 339402 700272 339408 700324
rect 339460 700312 339466 700324
rect 348786 700312 348792 700324
rect 339460 700284 348792 700312
rect 339460 700272 339466 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 351822 700272 351828 700324
rect 351880 700312 351886 700324
rect 364978 700312 364984 700324
rect 351880 700284 364984 700312
rect 351880 700272 351886 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 365622 700272 365628 700324
rect 365680 700312 365686 700324
rect 381170 700312 381176 700324
rect 365680 700284 381176 700312
rect 365680 700272 365686 700284
rect 381170 700272 381176 700284
rect 381228 700272 381234 700324
rect 390462 700272 390468 700324
rect 390520 700312 390526 700324
rect 413646 700312 413652 700324
rect 390520 700284 413652 700312
rect 390520 700272 390526 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 429102 700272 429108 700324
rect 429160 700312 429166 700324
rect 462314 700312 462320 700324
rect 429160 700284 462320 700312
rect 429160 700272 429166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 466362 700272 466368 700324
rect 466420 700312 466426 700324
rect 510982 700312 510988 700324
rect 466420 700284 510988 700312
rect 466420 700272 466426 700284
rect 510982 700272 510988 700284
rect 511040 700272 511046 700324
rect 517422 700272 517428 700324
rect 517480 700312 517486 700324
rect 575842 700312 575848 700324
rect 517480 700284 575848 700312
rect 517480 700272 517486 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 56778 700136 56784 700188
rect 56836 700176 56842 700188
rect 57882 700176 57888 700188
rect 56836 700148 57888 700176
rect 56836 700136 56842 700148
rect 57882 700136 57888 700148
rect 57940 700136 57946 700188
rect 186498 700136 186504 700188
rect 186556 700176 186562 700188
rect 187602 700176 187608 700188
rect 186556 700148 187608 700176
rect 186556 700136 186562 700148
rect 187602 700136 187608 700148
rect 187660 700136 187666 700188
rect 251450 700068 251456 700120
rect 251508 700108 251514 700120
rect 252462 700108 252468 700120
rect 251508 700080 252468 700108
rect 251508 700068 251514 700080
rect 252462 700068 252468 700080
rect 252520 700068 252526 700120
rect 283834 700068 283840 700120
rect 283892 700108 283898 700120
rect 284938 700108 284944 700120
rect 283892 700080 284944 700108
rect 283892 700068 283898 700080
rect 284938 700068 284944 700080
rect 284996 700068 285002 700120
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 314562 699660 314568 699712
rect 314620 699700 314626 699712
rect 316310 699700 316316 699712
rect 314620 699672 316316 699700
rect 314620 699660 314626 699672
rect 316310 699660 316316 699672
rect 316368 699660 316374 699712
rect 327718 699660 327724 699712
rect 327776 699700 327782 699712
rect 332502 699700 332508 699712
rect 327776 699672 332508 699700
rect 327776 699660 327782 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 519538 696940 519544 696992
rect 519596 696980 519602 696992
rect 580166 696980 580172 696992
rect 519596 696952 580172 696980
rect 519596 696940 519602 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 519630 683136 519636 683188
rect 519688 683176 519694 683188
rect 580166 683176 580172 683188
rect 519688 683148 580172 683176
rect 519688 683136 519694 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 519722 670692 519728 670744
rect 519780 670732 519786 670744
rect 580166 670732 580172 670744
rect 519780 670704 580172 670732
rect 519780 670692 519786 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 519814 656888 519820 656940
rect 519872 656928 519878 656940
rect 580166 656928 580172 656940
rect 519872 656900 580172 656928
rect 519872 656888 519878 656900
rect 580166 656888 580172 656900
rect 580224 656888 580230 656940
rect 519906 643084 519912 643136
rect 519964 643124 519970 643136
rect 580166 643124 580172 643136
rect 519964 643096 580172 643124
rect 519964 643084 519970 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 284938 643016 284944 643068
rect 284996 643056 285002 643068
rect 288158 643056 288164 643068
rect 284996 643028 288164 643056
rect 284996 643016 285002 643028
rect 288158 643016 288164 643028
rect 288216 643016 288222 643068
rect 57882 642540 57888 642592
rect 57940 642580 57946 642592
rect 110138 642580 110144 642592
rect 57940 642552 110144 642580
rect 57940 642540 57946 642552
rect 110138 642540 110144 642552
rect 110196 642540 110202 642592
rect 122742 642540 122748 642592
rect 122800 642580 122806 642592
rect 161014 642580 161020 642592
rect 122800 642552 161020 642580
rect 122800 642540 122806 642552
rect 161014 642540 161020 642552
rect 161072 642540 161078 642592
rect 440878 642540 440884 642592
rect 440936 642580 440942 642592
rect 441522 642580 441528 642592
rect 440936 642552 441528 642580
rect 440936 642540 440942 642552
rect 441522 642540 441528 642552
rect 441580 642540 441586 642592
rect 41322 642472 41328 642524
rect 41380 642512 41386 642524
rect 97350 642512 97356 642524
rect 41380 642484 97356 642512
rect 41380 642472 41386 642484
rect 97350 642472 97356 642484
rect 97408 642472 97414 642524
rect 106182 642472 106188 642524
rect 106240 642512 106246 642524
rect 148226 642512 148232 642524
rect 106240 642484 148232 642512
rect 106240 642472 106246 642484
rect 148226 642472 148232 642484
rect 148284 642472 148290 642524
rect 171042 642472 171048 642524
rect 171100 642512 171106 642524
rect 199102 642512 199108 642524
rect 171100 642484 199108 642512
rect 171100 642472 171106 642484
rect 199102 642472 199108 642484
rect 199160 642472 199166 642524
rect 24762 642404 24768 642456
rect 24820 642444 24826 642456
rect 84654 642444 84660 642456
rect 24820 642416 84660 642444
rect 24820 642404 24826 642416
rect 84654 642404 84660 642416
rect 84712 642404 84718 642456
rect 89622 642404 89628 642456
rect 89680 642444 89686 642456
rect 135530 642444 135536 642456
rect 89680 642416 135536 642444
rect 89680 642404 89686 642416
rect 135530 642404 135536 642416
rect 135588 642404 135594 642456
rect 154482 642404 154488 642456
rect 154540 642444 154546 642456
rect 186406 642444 186412 642456
rect 154540 642416 186412 642444
rect 154540 642404 154546 642416
rect 186406 642404 186412 642416
rect 186464 642404 186470 642456
rect 202782 642404 202788 642456
rect 202840 642444 202846 642456
rect 224586 642444 224592 642456
rect 202840 642416 224592 642444
rect 202840 642404 202846 642416
rect 224586 642404 224592 642416
rect 224644 642404 224650 642456
rect 235902 642404 235908 642456
rect 235960 642444 235966 642456
rect 249978 642444 249984 642456
rect 235960 642416 249984 642444
rect 235960 642404 235966 642416
rect 249978 642404 249984 642416
rect 250036 642404 250042 642456
rect 8202 642336 8208 642388
rect 8260 642376 8266 642388
rect 72786 642376 72792 642388
rect 8260 642348 72792 642376
rect 8260 642336 8266 642348
rect 72786 642336 72792 642348
rect 72844 642336 72850 642388
rect 73062 642336 73068 642388
rect 73120 642376 73126 642388
rect 122834 642376 122840 642388
rect 73120 642348 122840 642376
rect 73120 642336 73126 642348
rect 122834 642336 122840 642348
rect 122892 642336 122898 642388
rect 137922 642336 137928 642388
rect 137980 642376 137986 642388
rect 173710 642376 173716 642388
rect 137980 642348 173716 642376
rect 137980 642336 137986 642348
rect 173710 642336 173716 642348
rect 173768 642336 173774 642388
rect 187602 642336 187608 642388
rect 187660 642376 187666 642388
rect 211890 642376 211896 642388
rect 187660 642348 211896 642376
rect 187660 642336 187666 642348
rect 211890 642336 211896 642348
rect 211948 642336 211954 642388
rect 219342 642336 219348 642388
rect 219400 642376 219406 642388
rect 237282 642376 237288 642388
rect 219400 642348 237288 642376
rect 219400 642336 219406 642348
rect 237282 642336 237288 642348
rect 237340 642336 237346 642388
rect 252462 642336 252468 642388
rect 252520 642376 252526 642388
rect 262766 642376 262772 642388
rect 252520 642348 262772 642376
rect 252520 642336 252526 642348
rect 262766 642336 262772 642348
rect 262824 642336 262830 642388
rect 267642 642336 267648 642388
rect 267700 642376 267706 642388
rect 275462 642376 275468 642388
rect 267700 642348 275468 642376
rect 267700 642336 267706 642348
rect 275462 642336 275468 642348
rect 275520 642336 275526 642388
rect 313642 641724 313648 641776
rect 313700 641764 313706 641776
rect 314562 641764 314568 641776
rect 313700 641736 314568 641764
rect 313700 641724 313706 641736
rect 314562 641724 314568 641736
rect 314620 641724 314626 641776
rect 326338 641724 326344 641776
rect 326396 641764 326402 641776
rect 327718 641764 327724 641776
rect 326396 641736 327724 641764
rect 326396 641724 326402 641736
rect 327718 641724 327724 641736
rect 327776 641724 327782 641776
rect 364518 641724 364524 641776
rect 364576 641764 364582 641776
rect 365622 641764 365628 641776
rect 364576 641736 365628 641764
rect 364576 641724 364582 641736
rect 365622 641724 365628 641736
rect 365680 641724 365686 641776
rect 377214 641724 377220 641776
rect 377272 641764 377278 641776
rect 378042 641764 378048 641776
rect 377272 641736 378048 641764
rect 377272 641724 377278 641736
rect 378042 641724 378048 641736
rect 378100 641724 378106 641776
rect 390002 641724 390008 641776
rect 390060 641764 390066 641776
rect 390462 641764 390468 641776
rect 390060 641736 390468 641764
rect 390060 641724 390066 641736
rect 390462 641724 390468 641736
rect 390520 641724 390526 641776
rect 415394 641724 415400 641776
rect 415452 641764 415458 641776
rect 416682 641764 416688 641776
rect 415452 641736 416688 641764
rect 415452 641724 415458 641736
rect 416682 641724 416688 641736
rect 416740 641724 416746 641776
rect 428090 641724 428096 641776
rect 428148 641764 428154 641776
rect 429102 641764 429108 641776
rect 428148 641736 429108 641764
rect 428148 641724 428154 641736
rect 429102 641724 429108 641736
rect 429160 641724 429166 641776
rect 478966 641724 478972 641776
rect 479024 641764 479030 641776
rect 480162 641764 480168 641776
rect 479024 641736 480168 641764
rect 479024 641724 479030 641736
rect 480162 641724 480168 641736
rect 480220 641724 480226 641776
rect 491754 641724 491760 641776
rect 491812 641764 491818 641776
rect 492582 641764 492588 641776
rect 491812 641736 492588 641764
rect 491812 641724 491818 641736
rect 492582 641724 492588 641736
rect 492640 641724 492646 641776
rect 504450 641724 504456 641776
rect 504508 641764 504514 641776
rect 505002 641764 505008 641776
rect 504508 641736 505008 641764
rect 504508 641724 504514 641736
rect 505002 641724 505008 641736
rect 505060 641724 505066 641776
rect 516502 641724 516508 641776
rect 516560 641764 516566 641776
rect 517422 641764 517428 641776
rect 516560 641736 517428 641764
rect 516560 641724 516566 641736
rect 517422 641724 517428 641736
rect 517480 641724 517486 641776
rect 3418 637508 3424 637560
rect 3476 637548 3482 637560
rect 69014 637548 69020 637560
rect 3476 637520 69020 637548
rect 3476 637508 3482 637520
rect 69014 637508 69020 637520
rect 69072 637508 69078 637560
rect 519538 630640 519544 630692
rect 519596 630680 519602 630692
rect 580166 630680 580172 630692
rect 519596 630652 580172 630680
rect 519596 630640 519602 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 626492 3516 626544
rect 3568 626532 3574 626544
rect 69014 626532 69020 626544
rect 3568 626504 69020 626532
rect 3568 626492 3574 626504
rect 69014 626492 69020 626504
rect 69072 626492 69078 626544
rect 519630 616836 519636 616888
rect 519688 616876 519694 616888
rect 580166 616876 580172 616888
rect 519688 616848 580172 616876
rect 519688 616836 519694 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3602 615408 3608 615460
rect 3660 615448 3666 615460
rect 69014 615448 69020 615460
rect 3660 615420 69020 615448
rect 3660 615408 3666 615420
rect 69014 615408 69020 615420
rect 69072 615408 69078 615460
rect 3694 605752 3700 605804
rect 3752 605792 3758 605804
rect 69014 605792 69020 605804
rect 3752 605764 69020 605792
rect 3752 605752 3758 605764
rect 69014 605752 69020 605764
rect 69072 605752 69078 605804
rect 519722 603100 519728 603152
rect 519780 603140 519786 603152
rect 580166 603140 580172 603152
rect 519780 603112 580172 603140
rect 519780 603100 519786 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 3786 594736 3792 594788
rect 3844 594776 3850 594788
rect 69014 594776 69020 594788
rect 3844 594748 69020 594776
rect 3844 594736 3850 594748
rect 69014 594736 69020 594748
rect 69072 594736 69078 594788
rect 519814 590656 519820 590708
rect 519872 590696 519878 590708
rect 579798 590696 579804 590708
rect 519872 590668 579804 590696
rect 519872 590656 519878 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3418 583652 3424 583704
rect 3476 583692 3482 583704
rect 69014 583692 69020 583704
rect 3476 583664 69020 583692
rect 3476 583652 3482 583664
rect 69014 583652 69020 583664
rect 69072 583652 69078 583704
rect 519538 576852 519544 576904
rect 519596 576892 519602 576904
rect 580166 576892 580172 576904
rect 519596 576864 580172 576892
rect 519596 576852 519602 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3510 572636 3516 572688
rect 3568 572676 3574 572688
rect 69014 572676 69020 572688
rect 3568 572648 69020 572676
rect 3568 572636 3574 572648
rect 69014 572636 69020 572648
rect 69072 572636 69078 572688
rect 519630 563048 519636 563100
rect 519688 563088 519694 563100
rect 579798 563088 579804 563100
rect 519688 563060 579804 563088
rect 519688 563048 519694 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3602 561620 3608 561672
rect 3660 561660 3666 561672
rect 69014 561660 69020 561672
rect 3660 561632 69020 561660
rect 3660 561620 3666 561632
rect 69014 561620 69020 561632
rect 69072 561620 69078 561672
rect 519722 550604 519728 550656
rect 519780 550644 519786 550656
rect 580166 550644 580172 550656
rect 519780 550616 580172 550644
rect 519780 550604 519786 550616
rect 580166 550604 580172 550616
rect 580224 550604 580230 550656
rect 3694 550536 3700 550588
rect 3752 550576 3758 550588
rect 69014 550576 69020 550588
rect 3752 550548 69020 550576
rect 3752 550536 3758 550548
rect 69014 550536 69020 550548
rect 69072 550536 69078 550588
rect 3418 539520 3424 539572
rect 3476 539560 3482 539572
rect 69014 539560 69020 539572
rect 3476 539532 69020 539560
rect 3476 539520 3482 539532
rect 69014 539520 69020 539532
rect 69072 539520 69078 539572
rect 519814 536800 519820 536852
rect 519872 536840 519878 536852
rect 580166 536840 580172 536852
rect 519872 536812 580172 536840
rect 519872 536800 519878 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3510 528504 3516 528556
rect 3568 528544 3574 528556
rect 69014 528544 69020 528556
rect 3568 528516 69020 528544
rect 3568 528504 3574 528516
rect 69014 528504 69020 528516
rect 69072 528504 69078 528556
rect 519538 524424 519544 524476
rect 519596 524464 519602 524476
rect 580166 524464 580172 524476
rect 519596 524436 580172 524464
rect 519596 524424 519602 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3602 517420 3608 517472
rect 3660 517460 3666 517472
rect 69014 517460 69020 517472
rect 3660 517432 69020 517460
rect 3660 517420 3666 517432
rect 69014 517420 69020 517432
rect 69072 517420 69078 517472
rect 519630 510620 519636 510672
rect 519688 510660 519694 510672
rect 580166 510660 580172 510672
rect 519688 510632 580172 510660
rect 519688 510620 519694 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3694 507764 3700 507816
rect 3752 507804 3758 507816
rect 69014 507804 69020 507816
rect 3752 507776 69020 507804
rect 3752 507764 3758 507776
rect 69014 507764 69020 507776
rect 69072 507764 69078 507816
rect 519722 496816 519728 496868
rect 519780 496856 519786 496868
rect 580166 496856 580172 496868
rect 519780 496828 580172 496856
rect 519780 496816 519786 496828
rect 580166 496816 580172 496828
rect 580224 496816 580230 496868
rect 3418 496748 3424 496800
rect 3476 496788 3482 496800
rect 69014 496788 69020 496800
rect 3476 496760 69020 496788
rect 3476 496748 3482 496760
rect 69014 496748 69020 496760
rect 69072 496748 69078 496800
rect 3510 485732 3516 485784
rect 3568 485772 3574 485784
rect 69014 485772 69020 485784
rect 3568 485744 69020 485772
rect 3568 485732 3574 485744
rect 69014 485732 69020 485744
rect 69072 485732 69078 485784
rect 519538 484372 519544 484424
rect 519596 484412 519602 484424
rect 580166 484412 580172 484424
rect 519596 484384 580172 484412
rect 519596 484372 519602 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3602 474648 3608 474700
rect 3660 474688 3666 474700
rect 69014 474688 69020 474700
rect 3660 474660 69020 474688
rect 3660 474648 3666 474660
rect 69014 474648 69020 474660
rect 69072 474648 69078 474700
rect 519630 470568 519636 470620
rect 519688 470608 519694 470620
rect 579982 470608 579988 470620
rect 519688 470580 579988 470608
rect 519688 470568 519694 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3418 463632 3424 463684
rect 3476 463672 3482 463684
rect 69014 463672 69020 463684
rect 3476 463644 69020 463672
rect 3476 463632 3482 463644
rect 69014 463632 69020 463644
rect 69072 463632 69078 463684
rect 519538 456764 519544 456816
rect 519596 456804 519602 456816
rect 580166 456804 580172 456816
rect 519596 456776 580172 456804
rect 519596 456764 519602 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3510 452548 3516 452600
rect 3568 452588 3574 452600
rect 69014 452588 69020 452600
rect 3568 452560 69020 452588
rect 3568 452548 3574 452560
rect 69014 452548 69020 452560
rect 69072 452548 69078 452600
rect 519630 444388 519636 444440
rect 519688 444428 519694 444440
rect 580166 444428 580172 444440
rect 519688 444400 580172 444428
rect 519688 444388 519694 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 3602 441532 3608 441584
rect 3660 441572 3666 441584
rect 69014 441572 69020 441584
rect 3660 441544 69020 441572
rect 3660 441532 3666 441544
rect 69014 441532 69020 441544
rect 69072 441532 69078 441584
rect 519538 430584 519544 430636
rect 519596 430624 519602 430636
rect 580166 430624 580172 430636
rect 519596 430596 580172 430624
rect 519596 430584 519602 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 430516 3424 430568
rect 3476 430556 3482 430568
rect 69014 430556 69020 430568
rect 3476 430528 69020 430556
rect 3476 430516 3482 430528
rect 69014 430516 69020 430528
rect 69072 430516 69078 430568
rect 3510 419432 3516 419484
rect 3568 419472 3574 419484
rect 69014 419472 69020 419484
rect 3568 419444 69020 419472
rect 3568 419432 3574 419444
rect 69014 419432 69020 419444
rect 69072 419432 69078 419484
rect 519630 418140 519636 418192
rect 519688 418180 519694 418192
rect 580166 418180 580172 418192
rect 519688 418152 580172 418180
rect 519688 418140 519694 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3418 409776 3424 409828
rect 3476 409816 3482 409828
rect 69014 409816 69020 409828
rect 3476 409788 69020 409816
rect 3476 409776 3482 409788
rect 69014 409776 69020 409788
rect 69072 409776 69078 409828
rect 519538 404336 519544 404388
rect 519596 404376 519602 404388
rect 580166 404376 580172 404388
rect 519596 404348 580172 404376
rect 519596 404336 519602 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 398760 3516 398812
rect 3568 398800 3574 398812
rect 69014 398800 69020 398812
rect 3568 398772 69020 398800
rect 3568 398760 3574 398772
rect 69014 398760 69020 398772
rect 69072 398760 69078 398812
rect 519538 390532 519544 390584
rect 519596 390572 519602 390584
rect 580166 390572 580172 390584
rect 519596 390544 580172 390572
rect 519596 390532 519602 390544
rect 580166 390532 580172 390544
rect 580224 390532 580230 390584
rect 3418 387744 3424 387796
rect 3476 387784 3482 387796
rect 69014 387784 69020 387796
rect 3476 387756 69020 387784
rect 3476 387744 3482 387756
rect 69014 387744 69020 387756
rect 69072 387744 69078 387796
rect 519538 378156 519544 378208
rect 519596 378196 519602 378208
rect 580166 378196 580172 378208
rect 519596 378168 580172 378196
rect 519596 378156 519602 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 376660 3424 376712
rect 3476 376700 3482 376712
rect 69014 376700 69020 376712
rect 3476 376672 69020 376700
rect 3476 376660 3482 376672
rect 69014 376660 69020 376672
rect 69072 376660 69078 376712
rect 3418 365644 3424 365696
rect 3476 365684 3482 365696
rect 69014 365684 69020 365696
rect 3476 365656 69020 365684
rect 3476 365644 3482 365656
rect 69014 365644 69020 365656
rect 69072 365644 69078 365696
rect 519354 364352 519360 364404
rect 519412 364392 519418 364404
rect 580166 364392 580172 364404
rect 519412 364364 580172 364392
rect 519412 364352 519418 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 3418 354628 3424 354680
rect 3476 354668 3482 354680
rect 69014 354668 69020 354680
rect 3476 354640 69020 354668
rect 3476 354628 3482 354640
rect 69014 354628 69020 354640
rect 69072 354628 69078 354680
rect 519814 351908 519820 351960
rect 519872 351948 519878 351960
rect 580166 351948 580172 351960
rect 519872 351920 580172 351948
rect 519872 351908 519878 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3142 343544 3148 343596
rect 3200 343584 3206 343596
rect 69014 343584 69020 343596
rect 3200 343556 69020 343584
rect 3200 343544 3206 343556
rect 69014 343544 69020 343556
rect 69072 343544 69078 343596
rect 519998 338104 520004 338156
rect 520056 338144 520062 338156
rect 580166 338144 580172 338156
rect 520056 338116 580172 338144
rect 520056 338104 520062 338116
rect 580166 338104 580172 338116
rect 580224 338104 580230 338156
rect 3418 331848 3424 331900
rect 3476 331888 3482 331900
rect 69014 331888 69020 331900
rect 3476 331860 69020 331888
rect 3476 331848 3482 331860
rect 69014 331848 69020 331860
rect 69072 331848 69078 331900
rect 519354 325592 519360 325644
rect 519412 325632 519418 325644
rect 580166 325632 580172 325644
rect 519412 325604 580172 325632
rect 519412 325592 519418 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3418 320152 3424 320204
rect 3476 320192 3482 320204
rect 69014 320192 69020 320204
rect 3476 320164 69020 320192
rect 3476 320152 3482 320164
rect 69014 320152 69020 320164
rect 69072 320152 69078 320204
rect 520182 313216 520188 313268
rect 520240 313256 520246 313268
rect 580166 313256 580172 313268
rect 520240 313228 580172 313256
rect 520240 313216 520246 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3418 309136 3424 309188
rect 3476 309176 3482 309188
rect 69014 309176 69020 309188
rect 3476 309148 69020 309176
rect 3476 309136 3482 309148
rect 69014 309136 69020 309148
rect 69072 309136 69078 309188
rect 3418 299480 3424 299532
rect 3476 299520 3482 299532
rect 69014 299520 69020 299532
rect 3476 299492 69020 299520
rect 3476 299480 3482 299492
rect 69014 299480 69020 299492
rect 69072 299480 69078 299532
rect 519354 299412 519360 299464
rect 519412 299452 519418 299464
rect 580166 299452 580172 299464
rect 519412 299424 580172 299452
rect 519412 299412 519418 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3418 288396 3424 288448
rect 3476 288436 3482 288448
rect 69014 288436 69020 288448
rect 3476 288408 69020 288436
rect 3476 288396 3482 288408
rect 69014 288396 69020 288408
rect 69072 288396 69078 288448
rect 519538 285608 519544 285660
rect 519596 285648 519602 285660
rect 580166 285648 580172 285660
rect 519596 285620 580172 285648
rect 519596 285608 519602 285620
rect 580166 285608 580172 285620
rect 580224 285608 580230 285660
rect 3510 277380 3516 277432
rect 3568 277420 3574 277432
rect 69014 277420 69020 277432
rect 3568 277392 69020 277420
rect 3568 277380 3574 277392
rect 69014 277380 69020 277392
rect 69072 277380 69078 277432
rect 519538 273164 519544 273216
rect 519596 273204 519602 273216
rect 580166 273204 580172 273216
rect 519596 273176 580172 273204
rect 519596 273164 519602 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3418 266364 3424 266416
rect 3476 266404 3482 266416
rect 69014 266404 69020 266416
rect 3476 266376 69020 266404
rect 3476 266364 3482 266376
rect 69014 266364 69020 266376
rect 69072 266364 69078 266416
rect 519538 259360 519544 259412
rect 519596 259400 519602 259412
rect 580166 259400 580172 259412
rect 519596 259372 580172 259400
rect 519596 259360 519602 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3510 255280 3516 255332
rect 3568 255320 3574 255332
rect 69014 255320 69020 255332
rect 3568 255292 69020 255320
rect 3568 255280 3574 255292
rect 69014 255280 69020 255292
rect 69072 255280 69078 255332
rect 519630 245556 519636 245608
rect 519688 245596 519694 245608
rect 580166 245596 580172 245608
rect 519688 245568 580172 245596
rect 519688 245556 519694 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3418 244264 3424 244316
rect 3476 244304 3482 244316
rect 69014 244304 69020 244316
rect 3476 244276 69020 244304
rect 3476 244264 3482 244276
rect 69014 244264 69020 244276
rect 69072 244264 69078 244316
rect 3510 233248 3516 233300
rect 3568 233288 3574 233300
rect 69014 233288 69020 233300
rect 3568 233260 69020 233288
rect 3568 233248 3574 233260
rect 69014 233248 69020 233260
rect 69072 233248 69078 233300
rect 519538 233180 519544 233232
rect 519596 233220 519602 233232
rect 579982 233220 579988 233232
rect 519596 233192 579988 233220
rect 519596 233180 519602 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3418 222164 3424 222216
rect 3476 222204 3482 222216
rect 69014 222204 69020 222216
rect 3476 222176 69020 222204
rect 3476 222164 3482 222176
rect 69014 222164 69020 222176
rect 69072 222164 69078 222216
rect 519630 219376 519636 219428
rect 519688 219416 519694 219428
rect 580166 219416 580172 219428
rect 519688 219388 580172 219416
rect 519688 219376 519694 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3602 211148 3608 211200
rect 3660 211188 3666 211200
rect 69014 211188 69020 211200
rect 3660 211160 69020 211188
rect 3660 211148 3666 211160
rect 69014 211148 69020 211160
rect 69072 211148 69078 211200
rect 519538 206932 519544 206984
rect 519596 206972 519602 206984
rect 579798 206972 579804 206984
rect 519596 206944 579804 206972
rect 519596 206932 519602 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3510 201492 3516 201544
rect 3568 201532 3574 201544
rect 69014 201532 69020 201544
rect 3568 201504 69020 201532
rect 3568 201492 3574 201504
rect 69014 201492 69020 201504
rect 69072 201492 69078 201544
rect 519722 193128 519728 193180
rect 519780 193168 519786 193180
rect 580166 193168 580172 193180
rect 519780 193140 580172 193168
rect 519780 193128 519786 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3418 190476 3424 190528
rect 3476 190516 3482 190528
rect 69014 190516 69020 190528
rect 3476 190488 69020 190516
rect 3476 190476 3482 190488
rect 69014 190476 69020 190488
rect 69072 190476 69078 190528
rect 3602 179392 3608 179444
rect 3660 179432 3666 179444
rect 69014 179432 69020 179444
rect 3660 179404 69020 179432
rect 3660 179392 3666 179404
rect 69014 179392 69020 179404
rect 69072 179392 69078 179444
rect 519630 179324 519636 179376
rect 519688 179364 519694 179376
rect 580166 179364 580172 179376
rect 519688 179336 580172 179364
rect 519688 179324 519694 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 3510 168376 3516 168428
rect 3568 168416 3574 168428
rect 69014 168416 69020 168428
rect 3568 168388 69020 168416
rect 3568 168376 3574 168388
rect 69014 168376 69020 168388
rect 69072 168376 69078 168428
rect 519538 166948 519544 167000
rect 519596 166988 519602 167000
rect 580166 166988 580172 167000
rect 519596 166960 580172 166988
rect 519596 166948 519602 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3418 157360 3424 157412
rect 3476 157400 3482 157412
rect 69014 157400 69020 157412
rect 3476 157372 69020 157400
rect 3476 157360 3482 157372
rect 69014 157360 69020 157372
rect 69072 157360 69078 157412
rect 519722 153144 519728 153196
rect 519780 153184 519786 153196
rect 580166 153184 580172 153196
rect 519780 153156 580172 153184
rect 519780 153144 519786 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3694 146276 3700 146328
rect 3752 146316 3758 146328
rect 69014 146316 69020 146328
rect 3752 146288 69020 146316
rect 3752 146276 3758 146288
rect 69014 146276 69020 146288
rect 69072 146276 69078 146328
rect 519630 139340 519636 139392
rect 519688 139380 519694 139392
rect 580166 139380 580172 139392
rect 519688 139352 580172 139380
rect 519688 139340 519694 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3602 135260 3608 135312
rect 3660 135300 3666 135312
rect 69014 135300 69020 135312
rect 3660 135272 69020 135300
rect 3660 135260 3666 135272
rect 69014 135260 69020 135272
rect 69072 135260 69078 135312
rect 519538 126896 519544 126948
rect 519596 126936 519602 126948
rect 580166 126936 580172 126948
rect 519596 126908 580172 126936
rect 519596 126896 519602 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3510 124176 3516 124228
rect 3568 124216 3574 124228
rect 69014 124216 69020 124228
rect 3568 124188 69020 124216
rect 3568 124176 3574 124188
rect 69014 124176 69020 124188
rect 69072 124176 69078 124228
rect 3418 113160 3424 113212
rect 3476 113200 3482 113212
rect 69014 113200 69020 113212
rect 3476 113172 69020 113200
rect 3476 113160 3482 113172
rect 69014 113160 69020 113172
rect 69072 113160 69078 113212
rect 519814 113092 519820 113144
rect 519872 113132 519878 113144
rect 579798 113132 579804 113144
rect 519872 113104 579804 113132
rect 519872 113092 519878 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3786 103504 3792 103556
rect 3844 103544 3850 103556
rect 69014 103544 69020 103556
rect 3844 103516 69020 103544
rect 3844 103504 3850 103516
rect 69014 103504 69020 103516
rect 69072 103504 69078 103556
rect 519722 100648 519728 100700
rect 519780 100688 519786 100700
rect 580166 100688 580172 100700
rect 519780 100660 580172 100688
rect 519780 100648 519786 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3694 92488 3700 92540
rect 3752 92528 3758 92540
rect 69014 92528 69020 92540
rect 3752 92500 69020 92528
rect 3752 92488 3758 92500
rect 69014 92488 69020 92500
rect 69072 92488 69078 92540
rect 519630 86912 519636 86964
rect 519688 86952 519694 86964
rect 580166 86952 580172 86964
rect 519688 86924 580172 86952
rect 519688 86912 519694 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3602 81404 3608 81456
rect 3660 81444 3666 81456
rect 69014 81444 69020 81456
rect 3660 81416 69020 81444
rect 3660 81404 3666 81416
rect 69014 81404 69020 81416
rect 69072 81404 69078 81456
rect 519538 73108 519544 73160
rect 519596 73148 519602 73160
rect 580166 73148 580172 73160
rect 519596 73120 580172 73148
rect 519596 73108 519602 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 70388 3516 70440
rect 3568 70428 3574 70440
rect 69014 70428 69020 70440
rect 3568 70400 69020 70428
rect 3568 70388 3574 70400
rect 69014 70388 69020 70400
rect 69072 70388 69078 70440
rect 519906 60664 519912 60716
rect 519964 60704 519970 60716
rect 580166 60704 580172 60716
rect 519964 60676 580172 60704
rect 519964 60664 519970 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 303614 59848 303620 59900
rect 303672 59888 303678 59900
rect 304928 59888 304934 59900
rect 303672 59860 304934 59888
rect 303672 59848 303678 59860
rect 304928 59848 304934 59860
rect 304986 59848 304992 59900
rect 86954 59780 86960 59832
rect 87012 59820 87018 59832
rect 88208 59820 88214 59832
rect 87012 59792 88214 59820
rect 87012 59780 87018 59792
rect 88208 59780 88214 59792
rect 88266 59780 88272 59832
rect 89806 59780 89812 59832
rect 89864 59820 89870 59832
rect 90928 59820 90934 59832
rect 89864 59792 90934 59820
rect 89864 59780 89870 59792
rect 90928 59780 90934 59792
rect 90986 59780 90992 59832
rect 110414 59780 110420 59832
rect 110472 59820 110478 59832
rect 111688 59820 111694 59832
rect 110472 59792 111694 59820
rect 110472 59780 110478 59792
rect 111688 59780 111694 59792
rect 111746 59780 111752 59832
rect 133966 59780 133972 59832
rect 134024 59820 134030 59832
rect 135168 59820 135174 59832
rect 134024 59792 135174 59820
rect 134024 59780 134030 59792
rect 135168 59780 135174 59792
rect 135226 59780 135232 59832
rect 136634 59780 136640 59832
rect 136692 59820 136698 59832
rect 137868 59820 137874 59832
rect 136692 59792 137874 59820
rect 136692 59780 136698 59792
rect 137868 59780 137874 59792
rect 137926 59780 137932 59832
rect 139394 59780 139400 59832
rect 139452 59820 139458 59832
rect 140588 59820 140594 59832
rect 139452 59792 140594 59820
rect 139452 59780 139458 59792
rect 140588 59780 140594 59792
rect 140646 59780 140652 59832
rect 142154 59780 142160 59832
rect 142212 59820 142218 59832
rect 143288 59820 143294 59832
rect 142212 59792 143294 59820
rect 142212 59780 142218 59792
rect 143288 59780 143294 59792
rect 143346 59780 143352 59832
rect 150434 59780 150440 59832
rect 150492 59820 150498 59832
rect 151428 59820 151434 59832
rect 150492 59792 151434 59820
rect 150492 59780 150498 59792
rect 151428 59780 151434 59792
rect 151486 59780 151492 59832
rect 157334 59780 157340 59832
rect 157392 59820 157398 59832
rect 158648 59820 158654 59832
rect 157392 59792 158654 59820
rect 157392 59780 157398 59792
rect 158648 59780 158654 59792
rect 158706 59780 158712 59832
rect 160186 59780 160192 59832
rect 160244 59820 160250 59832
rect 161348 59820 161354 59832
rect 160244 59792 161354 59820
rect 160244 59780 160250 59792
rect 161348 59780 161354 59792
rect 161406 59780 161412 59832
rect 162946 59780 162952 59832
rect 163004 59820 163010 59832
rect 164068 59820 164074 59832
rect 163004 59792 164074 59820
rect 163004 59780 163010 59792
rect 164068 59780 164074 59792
rect 164126 59780 164132 59832
rect 168374 59780 168380 59832
rect 168432 59820 168438 59832
rect 169488 59820 169494 59832
rect 168432 59792 169494 59820
rect 168432 59780 168438 59792
rect 169488 59780 169494 59792
rect 169546 59780 169552 59832
rect 173894 59780 173900 59832
rect 173952 59820 173958 59832
rect 174908 59820 174914 59832
rect 173952 59792 174914 59820
rect 173952 59780 173958 59792
rect 174908 59780 174914 59792
rect 174966 59780 174972 59832
rect 291194 59780 291200 59832
rect 291252 59820 291258 59832
rect 292288 59820 292294 59832
rect 291252 59792 292294 59820
rect 291252 59780 291258 59792
rect 292288 59780 292294 59792
rect 292346 59780 292352 59832
rect 402974 59780 402980 59832
rect 403032 59820 403038 59832
rect 404268 59820 404274 59832
rect 403032 59792 404274 59820
rect 403032 59780 403038 59792
rect 404268 59780 404274 59792
rect 404326 59780 404332 59832
rect 405734 59780 405740 59832
rect 405792 59820 405798 59832
rect 406968 59820 406974 59832
rect 405792 59792 406974 59820
rect 405792 59780 405798 59792
rect 406968 59780 406974 59792
rect 407026 59780 407032 59832
rect 411254 59780 411260 59832
rect 411312 59820 411318 59832
rect 412388 59820 412394 59832
rect 411312 59792 412394 59820
rect 411312 59780 411318 59792
rect 412388 59780 412394 59792
rect 412446 59780 412452 59832
rect 414014 59780 414020 59832
rect 414072 59820 414078 59832
rect 415108 59820 415114 59832
rect 414072 59792 415114 59820
rect 414072 59780 414078 59792
rect 415108 59780 415114 59792
rect 415166 59780 415172 59832
rect 416774 59780 416780 59832
rect 416832 59820 416838 59832
rect 417808 59820 417814 59832
rect 416832 59792 417814 59820
rect 416832 59780 416838 59792
rect 417808 59780 417814 59792
rect 417866 59780 417872 59832
rect 419534 59780 419540 59832
rect 419592 59820 419598 59832
rect 420508 59820 420514 59832
rect 419592 59792 420514 59820
rect 419592 59780 419598 59792
rect 420508 59780 420514 59792
rect 420566 59780 420572 59832
rect 429194 59780 429200 59832
rect 429252 59820 429258 59832
rect 430448 59820 430454 59832
rect 429252 59792 430454 59820
rect 429252 59780 429258 59792
rect 430448 59780 430454 59792
rect 430506 59780 430512 59832
rect 431954 59780 431960 59832
rect 432012 59820 432018 59832
rect 433168 59820 433174 59832
rect 432012 59792 433174 59820
rect 432012 59780 432018 59792
rect 433168 59780 433174 59792
rect 433226 59780 433232 59832
rect 434714 59780 434720 59832
rect 434772 59820 434778 59832
rect 435868 59820 435874 59832
rect 434772 59792 435874 59820
rect 434772 59780 434778 59792
rect 435868 59780 435874 59792
rect 435926 59780 435932 59832
rect 442994 59780 443000 59832
rect 443052 59820 443058 59832
rect 443988 59820 443994 59832
rect 443052 59792 443994 59820
rect 443052 59780 443058 59792
rect 443988 59780 443994 59792
rect 444046 59780 444052 59832
rect 452654 59780 452660 59832
rect 452712 59820 452718 59832
rect 453928 59820 453934 59832
rect 452712 59792 453934 59820
rect 452712 59780 452718 59792
rect 453928 59780 453934 59792
rect 453986 59780 453992 59832
rect 463786 59780 463792 59832
rect 463844 59820 463850 59832
rect 464768 59820 464774 59832
rect 463844 59792 464774 59820
rect 463844 59780 463850 59792
rect 464768 59780 464774 59792
rect 464826 59780 464832 59832
rect 476206 59780 476212 59832
rect 476264 59820 476270 59832
rect 477408 59820 477414 59832
rect 476264 59792 477414 59820
rect 476264 59780 476270 59792
rect 477408 59780 477414 59792
rect 477466 59780 477472 59832
rect 3418 59372 3424 59424
rect 3476 59412 3482 59424
rect 69014 59412 69020 59424
rect 3476 59384 69020 59412
rect 3476 59372 3482 59384
rect 69014 59372 69020 59384
rect 69072 59372 69078 59424
rect 67545 57919 67603 57925
rect 67545 57885 67557 57919
rect 67591 57916 67603 57919
rect 72418 57916 72424 57928
rect 67591 57888 72424 57916
rect 67591 57885 67603 57888
rect 67545 57879 67603 57885
rect 72418 57876 72424 57888
rect 72476 57876 72482 57928
rect 72513 57919 72571 57925
rect 72513 57885 72525 57919
rect 72559 57916 72571 57919
rect 85482 57916 85488 57928
rect 72559 57888 85488 57916
rect 72559 57885 72571 57888
rect 72513 57879 72571 57885
rect 85482 57876 85488 57888
rect 85540 57876 85546 57928
rect 87598 57876 87604 57928
rect 87656 57916 87662 57928
rect 92474 57916 92480 57928
rect 87656 57888 92480 57916
rect 87656 57876 87662 57888
rect 92474 57876 92480 57888
rect 92532 57876 92538 57928
rect 100662 57876 100668 57928
rect 100720 57916 100726 57928
rect 106185 57919 106243 57925
rect 100720 57888 103514 57916
rect 100720 57876 100726 57888
rect 57238 57808 57244 57860
rect 57296 57848 57302 57860
rect 78306 57848 78312 57860
rect 57296 57820 78312 57848
rect 57296 57808 57302 57820
rect 78306 57808 78312 57820
rect 78364 57808 78370 57860
rect 88978 57808 88984 57860
rect 89036 57848 89042 57860
rect 91830 57848 91836 57860
rect 89036 57820 91836 57848
rect 89036 57808 89042 57820
rect 91830 57808 91836 57820
rect 91888 57808 91894 57860
rect 97258 57808 97264 57860
rect 97316 57848 97322 57860
rect 97902 57848 97908 57860
rect 97316 57820 97908 57848
rect 97316 57808 97322 57820
rect 97902 57808 97908 57820
rect 97960 57808 97966 57860
rect 98178 57808 98184 57860
rect 98236 57848 98242 57860
rect 99190 57848 99196 57860
rect 98236 57820 99196 57848
rect 98236 57808 98242 57820
rect 99190 57808 99196 57820
rect 99248 57808 99254 57860
rect 99926 57808 99932 57860
rect 99984 57848 99990 57860
rect 100570 57848 100576 57860
rect 99984 57820 100576 57848
rect 99984 57808 99990 57820
rect 100570 57808 100576 57820
rect 100628 57808 100634 57860
rect 100846 57808 100852 57860
rect 100904 57848 100910 57860
rect 102042 57848 102048 57860
rect 100904 57820 102048 57848
rect 100904 57808 100910 57820
rect 102042 57808 102048 57820
rect 102100 57808 102106 57860
rect 103486 57848 103514 57888
rect 106185 57885 106197 57919
rect 106231 57916 106243 57919
rect 109862 57916 109868 57928
rect 106231 57888 109868 57916
rect 106231 57885 106243 57888
rect 106185 57879 106243 57885
rect 109862 57876 109868 57888
rect 109920 57876 109926 57928
rect 213730 57876 213736 57928
rect 213788 57916 213794 57928
rect 305638 57916 305644 57928
rect 213788 57888 305644 57916
rect 213788 57876 213794 57888
rect 305638 57876 305644 57888
rect 305696 57876 305702 57928
rect 355502 57876 355508 57928
rect 355560 57916 355566 57928
rect 358078 57916 358084 57928
rect 355560 57888 358084 57916
rect 355560 57876 355566 57888
rect 358078 57876 358084 57888
rect 358136 57876 358142 57928
rect 363598 57876 363604 57928
rect 363656 57916 363662 57928
rect 364242 57916 364248 57928
rect 363656 57888 364248 57916
rect 363656 57876 363662 57888
rect 364242 57876 364248 57888
rect 364300 57876 364306 57928
rect 379882 57876 379888 57928
rect 379940 57916 379946 57928
rect 383565 57919 383623 57925
rect 383565 57916 383577 57919
rect 379940 57888 383577 57916
rect 379940 57876 379946 57888
rect 383565 57885 383577 57888
rect 383611 57885 383623 57919
rect 383565 57879 383623 57885
rect 392670 57876 392676 57928
rect 392728 57916 392734 57928
rect 402422 57916 402428 57928
rect 392728 57888 402428 57916
rect 392728 57876 392734 57888
rect 402422 57876 402428 57888
rect 402480 57876 402486 57928
rect 437658 57916 437664 57928
rect 431926 57888 437664 57916
rect 155034 57848 155040 57860
rect 103486 57820 155040 57848
rect 155034 57808 155040 57820
rect 155092 57808 155098 57860
rect 221826 57808 221832 57860
rect 221884 57848 221890 57860
rect 322198 57848 322204 57860
rect 221884 57820 322204 57848
rect 221884 57808 221890 57820
rect 322198 57808 322204 57820
rect 322256 57808 322262 57860
rect 353662 57808 353668 57860
rect 353720 57848 353726 57860
rect 378778 57848 378784 57860
rect 353720 57820 378784 57848
rect 353720 57808 353726 57820
rect 378778 57808 378784 57820
rect 378836 57808 378842 57860
rect 381538 57808 381544 57860
rect 381596 57848 381602 57860
rect 400674 57848 400680 57860
rect 381596 57820 400680 57848
rect 381596 57808 381602 57820
rect 400674 57808 400680 57820
rect 400732 57808 400738 57860
rect 431218 57808 431224 57860
rect 431276 57848 431282 57860
rect 431926 57848 431954 57888
rect 437658 57876 437664 57888
rect 437716 57876 437722 57928
rect 466362 57876 466368 57928
rect 466420 57916 466426 57928
rect 484578 57916 484584 57928
rect 466420 57888 484584 57916
rect 466420 57876 466426 57888
rect 484578 57876 484584 57888
rect 484636 57876 484642 57928
rect 431276 57820 431954 57848
rect 431276 57808 431282 57820
rect 436738 57808 436744 57860
rect 436796 57848 436802 57860
rect 438578 57848 438584 57860
rect 436796 57820 438584 57848
rect 436796 57808 436802 57820
rect 438578 57808 438584 57820
rect 438636 57808 438642 57860
rect 439498 57808 439504 57860
rect 439556 57848 439562 57860
rect 440418 57848 440424 57860
rect 439556 57820 440424 57848
rect 439556 57808 439562 57820
rect 440418 57808 440424 57820
rect 440476 57808 440482 57860
rect 441522 57808 441528 57860
rect 441580 57848 441586 57860
rect 478322 57848 478328 57860
rect 441580 57820 478328 57848
rect 441580 57808 441586 57820
rect 478322 57808 478328 57820
rect 478380 57808 478386 57860
rect 54478 57740 54484 57792
rect 54536 57780 54542 57792
rect 114370 57780 114376 57792
rect 54536 57752 114376 57780
rect 54536 57740 54542 57752
rect 114370 57740 114376 57752
rect 114428 57740 114434 57792
rect 225506 57740 225512 57792
rect 225564 57780 225570 57792
rect 340046 57780 340052 57792
rect 225564 57752 340052 57780
rect 225564 57740 225570 57752
rect 340046 57740 340052 57752
rect 340104 57740 340110 57792
rect 356422 57740 356428 57792
rect 356480 57780 356486 57792
rect 357250 57780 357256 57792
rect 356480 57752 357256 57780
rect 356480 57740 356486 57752
rect 357250 57740 357256 57752
rect 357308 57740 357314 57792
rect 358262 57740 358268 57792
rect 358320 57780 358326 57792
rect 358722 57780 358728 57792
rect 358320 57752 358728 57780
rect 358320 57740 358326 57752
rect 358722 57740 358728 57752
rect 358780 57740 358786 57792
rect 359090 57740 359096 57792
rect 359148 57780 359154 57792
rect 360102 57780 360108 57792
rect 359148 57752 360108 57780
rect 359148 57740 359154 57752
rect 360102 57740 360108 57752
rect 360160 57740 360166 57792
rect 360930 57740 360936 57792
rect 360988 57780 360994 57792
rect 361482 57780 361488 57792
rect 360988 57752 361488 57780
rect 360988 57740 360994 57752
rect 361482 57740 361488 57752
rect 361540 57740 361546 57792
rect 361850 57740 361856 57792
rect 361908 57780 361914 57792
rect 362862 57780 362868 57792
rect 361908 57752 362868 57780
rect 361908 57740 361914 57752
rect 362862 57740 362868 57752
rect 362920 57740 362926 57792
rect 363598 57740 363604 57792
rect 363656 57780 363662 57792
rect 451274 57780 451280 57792
rect 363656 57752 451280 57780
rect 363656 57740 363662 57752
rect 451274 57740 451280 57752
rect 451332 57740 451338 57792
rect 464617 57783 464675 57789
rect 464617 57749 464629 57783
rect 464663 57780 464675 57783
rect 468386 57780 468392 57792
rect 464663 57752 468392 57780
rect 464663 57749 464675 57752
rect 464617 57743 464675 57749
rect 468386 57740 468392 57752
rect 468444 57740 468450 57792
rect 468481 57783 468539 57789
rect 468481 57749 468493 57783
rect 468527 57780 468539 57783
rect 483750 57780 483756 57792
rect 468527 57752 483756 57780
rect 468527 57749 468539 57752
rect 468481 57743 468539 57749
rect 483750 57740 483756 57752
rect 483808 57740 483814 57792
rect 50338 57672 50344 57724
rect 50396 57712 50402 57724
rect 106185 57715 106243 57721
rect 106185 57712 106197 57715
rect 50396 57684 106197 57712
rect 50396 57672 50402 57684
rect 106185 57681 106197 57684
rect 106231 57681 106243 57715
rect 106185 57675 106243 57681
rect 106274 57672 106280 57724
rect 106332 57712 106338 57724
rect 107102 57712 107108 57724
rect 106332 57684 107108 57712
rect 106332 57672 106338 57684
rect 107102 57672 107108 57684
rect 107160 57672 107166 57724
rect 115198 57672 115204 57724
rect 115256 57712 115262 57724
rect 120718 57712 120724 57724
rect 115256 57684 120724 57712
rect 115256 57672 115262 57684
rect 120718 57672 120724 57684
rect 120776 57672 120782 57724
rect 155862 57672 155868 57724
rect 155920 57712 155926 57724
rect 290458 57712 290464 57724
rect 155920 57684 290464 57712
rect 155920 57672 155926 57684
rect 290458 57672 290464 57684
rect 290516 57672 290522 57724
rect 298738 57672 298744 57724
rect 298796 57712 298802 57724
rect 301409 57715 301467 57721
rect 298796 57684 301360 57712
rect 298796 57672 298802 57684
rect 53098 57604 53104 57656
rect 53156 57644 53162 57656
rect 113450 57644 113456 57656
rect 53156 57616 113456 57644
rect 53156 57604 53162 57616
rect 113450 57604 113456 57616
rect 113508 57604 113514 57656
rect 116578 57604 116584 57656
rect 116636 57644 116642 57656
rect 117958 57644 117964 57656
rect 116636 57616 117964 57644
rect 116636 57604 116642 57616
rect 117958 57604 117964 57616
rect 118016 57604 118022 57656
rect 123478 57604 123484 57656
rect 123536 57644 123542 57656
rect 124306 57644 124312 57656
rect 123536 57616 124312 57644
rect 123536 57604 123542 57616
rect 124306 57604 124312 57616
rect 124364 57604 124370 57656
rect 126238 57604 126244 57656
rect 126296 57644 126302 57656
rect 127066 57644 127072 57656
rect 126296 57616 127072 57644
rect 126296 57604 126302 57616
rect 127066 57604 127072 57616
rect 127124 57604 127130 57656
rect 129734 57604 129740 57656
rect 129792 57644 129798 57656
rect 130654 57644 130660 57656
rect 129792 57616 130660 57644
rect 129792 57604 129798 57616
rect 130654 57604 130660 57616
rect 130712 57604 130718 57656
rect 144178 57604 144184 57656
rect 144236 57644 144242 57656
rect 145098 57644 145104 57656
rect 144236 57616 145104 57644
rect 144236 57604 144242 57616
rect 145098 57604 145104 57616
rect 145156 57604 145162 57656
rect 153194 57604 153200 57656
rect 153252 57644 153258 57656
rect 154114 57644 154120 57656
rect 153252 57616 154120 57644
rect 153252 57604 153258 57616
rect 154114 57604 154120 57616
rect 154172 57604 154178 57656
rect 166258 57604 166264 57656
rect 166316 57644 166322 57656
rect 167638 57644 167644 57656
rect 166316 57616 167644 57644
rect 166316 57604 166322 57616
rect 167638 57604 167644 57616
rect 167696 57604 167702 57656
rect 185762 57604 185768 57656
rect 185820 57644 185826 57656
rect 186958 57644 186964 57656
rect 185820 57616 186964 57644
rect 185820 57604 185826 57616
rect 186958 57604 186964 57616
rect 187016 57604 187022 57656
rect 191190 57604 191196 57656
rect 191248 57644 191254 57656
rect 191742 57644 191748 57656
rect 191248 57616 191748 57644
rect 191248 57604 191254 57616
rect 191742 57604 191748 57616
rect 191800 57604 191806 57656
rect 192018 57604 192024 57656
rect 192076 57644 192082 57656
rect 193030 57644 193036 57656
rect 192076 57616 193036 57644
rect 192076 57604 192082 57616
rect 193030 57604 193036 57616
rect 193088 57604 193094 57656
rect 193858 57604 193864 57656
rect 193916 57644 193922 57656
rect 194502 57644 194508 57656
rect 193916 57616 194508 57644
rect 193916 57604 193922 57616
rect 194502 57604 194508 57616
rect 194560 57604 194566 57656
rect 194778 57604 194784 57656
rect 194836 57644 194842 57656
rect 195790 57644 195796 57656
rect 194836 57616 195796 57644
rect 194836 57604 194842 57616
rect 195790 57604 195796 57616
rect 195848 57604 195854 57656
rect 196618 57604 196624 57656
rect 196676 57644 196682 57656
rect 197262 57644 197268 57656
rect 196676 57616 197268 57644
rect 196676 57604 196682 57616
rect 197262 57604 197268 57616
rect 197320 57604 197326 57656
rect 197446 57604 197452 57656
rect 197504 57644 197510 57656
rect 198642 57644 198648 57656
rect 197504 57616 198648 57644
rect 197504 57604 197510 57616
rect 198642 57604 198648 57616
rect 198700 57604 198706 57656
rect 199286 57604 199292 57656
rect 199344 57644 199350 57656
rect 200022 57644 200028 57656
rect 199344 57616 200028 57644
rect 199344 57604 199350 57616
rect 200022 57604 200028 57616
rect 200080 57604 200086 57656
rect 200206 57604 200212 57656
rect 200264 57644 200270 57656
rect 201402 57644 201408 57656
rect 200264 57616 201408 57644
rect 200264 57604 200270 57616
rect 201402 57604 201408 57616
rect 201460 57604 201466 57656
rect 202046 57604 202052 57656
rect 202104 57644 202110 57656
rect 202782 57644 202788 57656
rect 202104 57616 202788 57644
rect 202104 57604 202110 57616
rect 202782 57604 202788 57616
rect 202840 57604 202846 57656
rect 202874 57604 202880 57656
rect 202932 57644 202938 57656
rect 204162 57644 204168 57656
rect 202932 57616 204168 57644
rect 202932 57604 202938 57616
rect 204162 57604 204168 57616
rect 204220 57604 204226 57656
rect 204714 57604 204720 57656
rect 204772 57644 204778 57656
rect 205542 57644 205548 57656
rect 204772 57616 205548 57644
rect 204772 57604 204778 57616
rect 205542 57604 205548 57616
rect 205600 57604 205606 57656
rect 205634 57604 205640 57656
rect 205692 57644 205698 57656
rect 206830 57644 206836 57656
rect 205692 57616 206836 57644
rect 205692 57604 205698 57616
rect 206830 57604 206836 57616
rect 206888 57604 206894 57656
rect 207382 57604 207388 57656
rect 207440 57644 207446 57656
rect 208302 57644 208308 57656
rect 207440 57616 208308 57644
rect 207440 57604 207446 57616
rect 208302 57604 208308 57616
rect 208360 57604 208366 57656
rect 209222 57604 209228 57656
rect 209280 57644 209286 57656
rect 209682 57644 209688 57656
rect 209280 57616 209688 57644
rect 209280 57604 209286 57616
rect 209682 57604 209688 57616
rect 209740 57604 209746 57656
rect 212810 57604 212816 57656
rect 212868 57644 212874 57656
rect 213822 57644 213828 57656
rect 212868 57616 213828 57644
rect 212868 57604 212874 57616
rect 213822 57604 213828 57616
rect 213880 57604 213886 57656
rect 214650 57604 214656 57656
rect 214708 57644 214714 57656
rect 215202 57644 215208 57656
rect 214708 57616 215208 57644
rect 214708 57604 214714 57616
rect 215202 57604 215208 57616
rect 215260 57604 215266 57656
rect 215570 57604 215576 57656
rect 215628 57644 215634 57656
rect 216490 57644 216496 57656
rect 215628 57616 216496 57644
rect 215628 57604 215634 57616
rect 216490 57604 216496 57616
rect 216548 57604 216554 57656
rect 217318 57604 217324 57656
rect 217376 57644 217382 57656
rect 217962 57644 217968 57656
rect 217376 57616 217968 57644
rect 217376 57604 217382 57616
rect 217962 57604 217968 57616
rect 218020 57604 218026 57656
rect 220078 57604 220084 57656
rect 220136 57644 220142 57656
rect 220722 57644 220728 57656
rect 220136 57616 220728 57644
rect 220136 57604 220142 57616
rect 220722 57604 220728 57616
rect 220780 57604 220786 57656
rect 222746 57604 222752 57656
rect 222804 57644 222810 57656
rect 223482 57644 223488 57656
rect 222804 57616 223488 57644
rect 222804 57604 222810 57616
rect 223482 57604 223488 57616
rect 223540 57604 223546 57656
rect 223666 57604 223672 57656
rect 223724 57644 223730 57656
rect 224770 57644 224776 57656
rect 223724 57616 224776 57644
rect 223724 57604 223730 57616
rect 224770 57604 224776 57616
rect 224828 57604 224834 57656
rect 226426 57604 226432 57656
rect 226484 57644 226490 57656
rect 227530 57644 227536 57656
rect 226484 57616 227536 57644
rect 226484 57604 226490 57616
rect 227530 57604 227536 57616
rect 227588 57604 227594 57656
rect 228174 57604 228180 57656
rect 228232 57644 228238 57656
rect 229002 57644 229008 57656
rect 228232 57616 229008 57644
rect 228232 57604 228238 57616
rect 229002 57604 229008 57616
rect 229060 57604 229066 57656
rect 229094 57604 229100 57656
rect 229152 57644 229158 57656
rect 230290 57644 230296 57656
rect 229152 57616 230296 57644
rect 229152 57604 229158 57616
rect 230290 57604 230296 57616
rect 230348 57604 230354 57656
rect 230934 57604 230940 57656
rect 230992 57644 230998 57656
rect 231670 57644 231676 57656
rect 230992 57616 231676 57644
rect 230992 57604 230998 57616
rect 231670 57604 231676 57616
rect 231728 57604 231734 57656
rect 232682 57604 232688 57656
rect 232740 57644 232746 57656
rect 233142 57644 233148 57656
rect 232740 57616 233148 57644
rect 232740 57604 232746 57616
rect 233142 57604 233148 57616
rect 233200 57604 233206 57656
rect 236362 57604 236368 57656
rect 236420 57644 236426 57656
rect 238018 57644 238024 57656
rect 236420 57616 238024 57644
rect 236420 57604 236426 57616
rect 238018 57604 238024 57616
rect 238076 57604 238082 57656
rect 238205 57647 238263 57653
rect 238205 57613 238217 57647
rect 238251 57644 238263 57647
rect 301225 57647 301283 57653
rect 301225 57644 301237 57647
rect 238251 57616 301237 57644
rect 238251 57613 238263 57616
rect 238205 57607 238263 57613
rect 301225 57613 301237 57616
rect 301271 57613 301283 57647
rect 301225 57607 301283 57613
rect 11698 57536 11704 57588
rect 11756 57576 11762 57588
rect 67545 57579 67603 57585
rect 67545 57576 67557 57579
rect 11756 57548 67557 57576
rect 11756 57536 11762 57548
rect 67545 57545 67557 57548
rect 67591 57545 67603 57579
rect 67545 57539 67603 57545
rect 71038 57536 71044 57588
rect 71096 57576 71102 57588
rect 73798 57576 73804 57588
rect 71096 57548 73804 57576
rect 71096 57536 71102 57548
rect 73798 57536 73804 57548
rect 73856 57536 73862 57588
rect 79318 57536 79324 57588
rect 79376 57576 79382 57588
rect 115934 57576 115940 57588
rect 79376 57548 115940 57576
rect 79376 57536 79382 57548
rect 115934 57536 115940 57548
rect 115992 57536 115998 57588
rect 124858 57536 124864 57588
rect 124916 57576 124922 57588
rect 127894 57576 127900 57588
rect 124916 57548 127900 57576
rect 124916 57536 124922 57548
rect 127894 57536 127900 57548
rect 127952 57536 127958 57588
rect 128998 57536 129004 57588
rect 129056 57576 129062 57588
rect 131574 57576 131580 57588
rect 129056 57548 131580 57576
rect 129056 57536 129062 57548
rect 131574 57536 131580 57548
rect 131632 57536 131638 57588
rect 148962 57536 148968 57588
rect 149020 57576 149026 57588
rect 288434 57576 288440 57588
rect 149020 57548 288440 57576
rect 149020 57536 149026 57548
rect 288434 57536 288440 57548
rect 288492 57536 288498 57588
rect 289078 57536 289084 57588
rect 289136 57576 289142 57588
rect 293954 57576 293960 57588
rect 289136 57548 293960 57576
rect 289136 57536 289142 57548
rect 293954 57536 293960 57548
rect 294012 57536 294018 57588
rect 299474 57536 299480 57588
rect 299532 57576 299538 57588
rect 300394 57576 300400 57588
rect 299532 57548 300400 57576
rect 299532 57536 299538 57548
rect 300394 57536 300400 57548
rect 300452 57536 300458 57588
rect 301332 57576 301360 57684
rect 301409 57681 301421 57715
rect 301455 57712 301467 57715
rect 301455 57684 306374 57712
rect 301455 57681 301467 57684
rect 301409 57675 301467 57681
rect 306346 57644 306374 57684
rect 306466 57672 306472 57724
rect 306524 57712 306530 57724
rect 307662 57712 307668 57724
rect 306524 57684 307668 57712
rect 306524 57672 306530 57684
rect 307662 57672 307668 57684
rect 307720 57672 307726 57724
rect 331858 57672 331864 57724
rect 331916 57712 331922 57724
rect 333790 57712 333796 57724
rect 331916 57684 333796 57712
rect 331916 57672 331922 57684
rect 333790 57672 333796 57684
rect 333848 57672 333854 57724
rect 343818 57672 343824 57724
rect 343876 57712 343882 57724
rect 344922 57712 344928 57724
rect 343876 57684 344928 57712
rect 343876 57672 343882 57684
rect 344922 57672 344928 57684
rect 344980 57672 344986 57724
rect 345566 57672 345572 57724
rect 345624 57712 345630 57724
rect 346302 57712 346308 57724
rect 345624 57684 346308 57712
rect 345624 57672 345630 57684
rect 346302 57672 346308 57684
rect 346360 57672 346366 57724
rect 346486 57672 346492 57724
rect 346544 57712 346550 57724
rect 347682 57712 347688 57724
rect 346544 57684 347688 57712
rect 346544 57672 346550 57684
rect 347682 57672 347688 57684
rect 347740 57672 347746 57724
rect 348326 57672 348332 57724
rect 348384 57712 348390 57724
rect 349062 57712 349068 57724
rect 348384 57684 349068 57712
rect 348384 57672 348390 57684
rect 349062 57672 349068 57684
rect 349120 57672 349126 57724
rect 349246 57672 349252 57724
rect 349304 57712 349310 57724
rect 350350 57712 350356 57724
rect 349304 57684 350356 57712
rect 349304 57672 349310 57684
rect 350350 57672 350356 57684
rect 350408 57672 350414 57724
rect 350994 57672 351000 57724
rect 351052 57712 351058 57724
rect 351822 57712 351828 57724
rect 351052 57684 351828 57712
rect 351052 57672 351058 57684
rect 351822 57672 351828 57684
rect 351880 57672 351886 57724
rect 351914 57672 351920 57724
rect 351972 57712 351978 57724
rect 353202 57712 353208 57724
rect 351972 57684 353208 57712
rect 351972 57672 351978 57684
rect 353202 57672 353208 57684
rect 353260 57672 353266 57724
rect 353938 57672 353944 57724
rect 353996 57712 354002 57724
rect 445754 57712 445760 57724
rect 353996 57684 445760 57712
rect 353996 57672 354002 57684
rect 445754 57672 445760 57684
rect 445812 57672 445818 57724
rect 458082 57672 458088 57724
rect 458140 57712 458146 57724
rect 482830 57712 482836 57724
rect 458140 57684 482836 57712
rect 458140 57672 458146 57684
rect 482830 57672 482836 57684
rect 482888 57672 482894 57724
rect 364429 57647 364487 57653
rect 364429 57644 364441 57647
rect 306346 57616 364441 57644
rect 364429 57613 364441 57616
rect 364475 57613 364487 57647
rect 364429 57607 364487 57613
rect 364518 57604 364524 57656
rect 364576 57644 364582 57656
rect 365530 57644 365536 57656
rect 364576 57616 365536 57644
rect 364576 57604 364582 57616
rect 365530 57604 365536 57616
rect 365588 57604 365594 57656
rect 366358 57604 366364 57656
rect 366416 57644 366422 57656
rect 367002 57644 367008 57656
rect 366416 57616 367008 57644
rect 366416 57604 366422 57616
rect 367002 57604 367008 57616
rect 367060 57604 367066 57656
rect 367278 57604 367284 57656
rect 367336 57644 367342 57656
rect 368382 57644 368388 57656
rect 367336 57616 368388 57644
rect 367336 57604 367342 57616
rect 368382 57604 368388 57616
rect 368440 57604 368446 57656
rect 369026 57604 369032 57656
rect 369084 57644 369090 57656
rect 369762 57644 369768 57656
rect 369084 57616 369768 57644
rect 369084 57604 369090 57616
rect 369762 57604 369768 57616
rect 369820 57604 369826 57656
rect 369946 57604 369952 57656
rect 370004 57644 370010 57656
rect 371142 57644 371148 57656
rect 370004 57616 371148 57644
rect 370004 57604 370010 57616
rect 371142 57604 371148 57616
rect 371200 57604 371206 57656
rect 371786 57604 371792 57656
rect 371844 57644 371850 57656
rect 372522 57644 372528 57656
rect 371844 57616 372528 57644
rect 371844 57604 371850 57616
rect 372522 57604 372528 57616
rect 372580 57604 372586 57656
rect 372706 57604 372712 57656
rect 372764 57644 372770 57656
rect 373902 57644 373908 57656
rect 372764 57616 373908 57644
rect 372764 57604 372770 57616
rect 373902 57604 373908 57616
rect 373960 57604 373966 57656
rect 374454 57604 374460 57656
rect 374512 57644 374518 57656
rect 375282 57644 375288 57656
rect 374512 57616 375288 57644
rect 374512 57604 374518 57616
rect 375282 57604 375288 57616
rect 375340 57604 375346 57656
rect 375374 57604 375380 57656
rect 375432 57644 375438 57656
rect 376570 57644 376576 57656
rect 375432 57616 376576 57644
rect 375432 57604 375438 57616
rect 376570 57604 376576 57616
rect 376628 57604 376634 57656
rect 377214 57604 377220 57656
rect 377272 57644 377278 57656
rect 377950 57644 377956 57656
rect 377272 57616 377956 57644
rect 377272 57604 377278 57616
rect 377950 57604 377956 57616
rect 378008 57604 378014 57656
rect 378962 57604 378968 57656
rect 379020 57644 379026 57656
rect 379422 57644 379428 57656
rect 379020 57616 379428 57644
rect 379020 57604 379026 57616
rect 379422 57604 379428 57616
rect 379480 57604 379486 57656
rect 381722 57604 381728 57656
rect 381780 57644 381786 57656
rect 382182 57644 382188 57656
rect 381780 57616 382188 57644
rect 381780 57604 381786 57616
rect 382182 57604 382188 57616
rect 382240 57604 382246 57656
rect 382642 57604 382648 57656
rect 382700 57644 382706 57656
rect 383470 57644 383476 57656
rect 382700 57616 383476 57644
rect 382700 57604 382706 57616
rect 383470 57604 383476 57616
rect 383528 57604 383534 57656
rect 383565 57647 383623 57653
rect 383565 57613 383577 57647
rect 383611 57644 383623 57647
rect 418798 57644 418804 57656
rect 383611 57616 418804 57644
rect 383611 57613 383623 57616
rect 383565 57607 383623 57613
rect 418798 57604 418804 57616
rect 418856 57604 418862 57656
rect 425054 57604 425060 57656
rect 425112 57644 425118 57656
rect 425882 57644 425888 57656
rect 425112 57616 425888 57644
rect 425112 57604 425118 57616
rect 425882 57604 425888 57616
rect 425940 57604 425946 57656
rect 430482 57604 430488 57656
rect 430540 57644 430546 57656
rect 430540 57616 471928 57644
rect 430540 57604 430546 57616
rect 317414 57576 317420 57588
rect 301332 57548 317420 57576
rect 317414 57536 317420 57548
rect 317472 57536 317478 57588
rect 322934 57536 322940 57588
rect 322992 57576 322998 57588
rect 323854 57576 323860 57588
rect 322992 57548 323860 57576
rect 322992 57536 322998 57548
rect 323854 57536 323860 57548
rect 323912 57536 323918 57588
rect 325694 57536 325700 57588
rect 325752 57576 325758 57588
rect 326614 57576 326620 57588
rect 325752 57548 326620 57576
rect 325752 57536 325758 57548
rect 326614 57536 326620 57548
rect 326672 57536 326678 57588
rect 329926 57536 329932 57588
rect 329984 57576 329990 57588
rect 331122 57576 331128 57588
rect 329984 57548 331128 57576
rect 329984 57536 329990 57548
rect 331122 57536 331128 57548
rect 331180 57536 331186 57588
rect 335354 57536 335360 57588
rect 335412 57576 335418 57588
rect 336550 57576 336556 57588
rect 335412 57548 336556 57576
rect 335412 57536 335418 57548
rect 336550 57536 336556 57548
rect 336608 57536 336614 57588
rect 337470 57536 337476 57588
rect 337528 57576 337534 57588
rect 338022 57576 338028 57588
rect 337528 57548 338028 57576
rect 337528 57536 337534 57548
rect 338022 57536 338028 57548
rect 338080 57536 338086 57588
rect 338390 57536 338396 57588
rect 338448 57576 338454 57588
rect 339310 57576 339316 57588
rect 338448 57548 339316 57576
rect 338448 57536 338454 57548
rect 339310 57536 339316 57548
rect 339368 57536 339374 57588
rect 340138 57536 340144 57588
rect 340196 57576 340202 57588
rect 340782 57576 340788 57588
rect 340196 57548 340788 57576
rect 340196 57536 340202 57548
rect 340782 57536 340788 57548
rect 340840 57536 340846 57588
rect 341058 57536 341064 57588
rect 341116 57576 341122 57588
rect 342070 57576 342076 57588
rect 341116 57548 342076 57576
rect 341116 57536 341122 57548
rect 342070 57536 342076 57548
rect 342128 57536 342134 57588
rect 342898 57536 342904 57588
rect 342956 57576 342962 57588
rect 343542 57576 343548 57588
rect 342956 57548 343548 57576
rect 342956 57536 342962 57548
rect 343542 57536 343548 57548
rect 343600 57536 343606 57588
rect 344005 57579 344063 57585
rect 344005 57545 344017 57579
rect 344051 57576 344063 57579
rect 444834 57576 444840 57588
rect 344051 57548 444840 57576
rect 344051 57545 344063 57548
rect 344005 57539 344063 57545
rect 444834 57536 444840 57548
rect 444892 57536 444898 57588
rect 448514 57536 448520 57588
rect 448572 57576 448578 57588
rect 449342 57576 449348 57588
rect 448572 57548 449348 57576
rect 448572 57536 448578 57548
rect 449342 57536 449348 57548
rect 449400 57536 449406 57588
rect 449437 57579 449495 57585
rect 449437 57545 449449 57579
rect 449483 57576 449495 57579
rect 471793 57579 471851 57585
rect 471793 57576 471805 57579
rect 449483 57548 471805 57576
rect 449483 57545 449495 57548
rect 449437 57539 449495 57545
rect 471793 57545 471805 57548
rect 471839 57545 471851 57579
rect 471900 57576 471928 57616
rect 471974 57604 471980 57656
rect 472032 57644 472038 57656
rect 472894 57644 472900 57656
rect 472032 57616 472900 57644
rect 472032 57604 472038 57616
rect 472894 57604 472900 57616
rect 472952 57604 472958 57656
rect 480162 57604 480168 57656
rect 480220 57644 480226 57656
rect 488258 57644 488264 57656
rect 480220 57616 488264 57644
rect 480220 57604 480226 57616
rect 488258 57604 488264 57616
rect 488316 57604 488322 57656
rect 491846 57604 491852 57656
rect 491904 57644 491910 57656
rect 492858 57644 492864 57656
rect 491904 57616 492864 57644
rect 491904 57604 491910 57616
rect 492858 57604 492864 57616
rect 492916 57604 492922 57656
rect 494606 57604 494612 57656
rect 494664 57644 494670 57656
rect 495342 57644 495348 57656
rect 494664 57616 495348 57644
rect 494664 57604 494670 57616
rect 495342 57604 495348 57616
rect 495400 57604 495406 57656
rect 495526 57604 495532 57656
rect 495584 57644 495590 57656
rect 496722 57644 496728 57656
rect 495584 57616 496728 57644
rect 495584 57604 495590 57616
rect 496722 57604 496728 57616
rect 496780 57604 496786 57656
rect 497274 57604 497280 57656
rect 497332 57644 497338 57656
rect 498102 57644 498108 57656
rect 497332 57616 498108 57644
rect 497332 57604 497338 57616
rect 498102 57604 498108 57616
rect 498160 57604 498166 57656
rect 498194 57604 498200 57656
rect 498252 57644 498258 57656
rect 499390 57644 499396 57656
rect 498252 57616 499396 57644
rect 498252 57604 498258 57616
rect 499390 57604 499396 57616
rect 499448 57604 499454 57656
rect 500034 57604 500040 57656
rect 500092 57644 500098 57656
rect 500770 57644 500776 57656
rect 500092 57616 500776 57644
rect 500092 57604 500098 57616
rect 500770 57604 500776 57616
rect 500828 57604 500834 57656
rect 501782 57604 501788 57656
rect 501840 57644 501846 57656
rect 502242 57644 502248 57656
rect 501840 57616 502248 57644
rect 501840 57604 501846 57616
rect 502242 57604 502248 57616
rect 502300 57604 502306 57656
rect 505462 57604 505468 57656
rect 505520 57644 505526 57656
rect 506382 57644 506388 57656
rect 505520 57616 506388 57644
rect 505520 57604 505526 57616
rect 506382 57604 506388 57616
rect 506440 57604 506446 57656
rect 507210 57604 507216 57656
rect 507268 57644 507274 57656
rect 507762 57644 507768 57656
rect 507268 57616 507768 57644
rect 507268 57604 507274 57616
rect 507762 57604 507768 57616
rect 507820 57604 507826 57656
rect 508130 57604 508136 57656
rect 508188 57644 508194 57656
rect 509050 57644 509056 57656
rect 508188 57616 509056 57644
rect 508188 57604 508194 57616
rect 509050 57604 509056 57616
rect 509108 57604 509114 57656
rect 509878 57604 509884 57656
rect 509936 57644 509942 57656
rect 510522 57644 510528 57656
rect 509936 57616 510528 57644
rect 509936 57604 509942 57616
rect 510522 57604 510528 57616
rect 510580 57604 510586 57656
rect 510798 57604 510804 57656
rect 510856 57644 510862 57656
rect 511810 57644 511816 57656
rect 510856 57616 511816 57644
rect 510856 57604 510862 57616
rect 511810 57604 511816 57616
rect 511868 57604 511874 57656
rect 513558 57604 513564 57656
rect 513616 57644 513622 57656
rect 514570 57644 514576 57656
rect 513616 57616 514576 57644
rect 513616 57604 513622 57616
rect 514570 57604 514576 57616
rect 514628 57604 514634 57656
rect 515306 57604 515312 57656
rect 515364 57644 515370 57656
rect 516042 57644 516048 57656
rect 515364 57616 516048 57644
rect 515364 57604 515370 57616
rect 516042 57604 516048 57616
rect 516100 57604 516106 57656
rect 516870 57604 516876 57656
rect 516928 57644 516934 57656
rect 517422 57644 517428 57656
rect 516928 57616 517428 57644
rect 516928 57604 516934 57616
rect 517422 57604 517428 57616
rect 517480 57604 517486 57656
rect 475562 57576 475568 57588
rect 471900 57548 475568 57576
rect 471793 57539 471851 57545
rect 475562 57536 475568 57548
rect 475620 57536 475626 57588
rect 482922 57536 482928 57588
rect 482980 57576 482986 57588
rect 489178 57576 489184 57588
rect 482980 57548 489184 57576
rect 482980 57536 482986 57548
rect 489178 57536 489184 57548
rect 489236 57536 489242 57588
rect 492766 57536 492772 57588
rect 492824 57576 492830 57588
rect 493870 57576 493876 57588
rect 492824 57548 493876 57576
rect 492824 57536 492830 57548
rect 493870 57536 493876 57548
rect 493928 57536 493934 57588
rect 516226 57536 516232 57588
rect 516284 57576 516290 57588
rect 517330 57576 517336 57588
rect 516284 57548 517336 57576
rect 516284 57536 516290 57548
rect 517330 57536 517336 57548
rect 517388 57536 517394 57588
rect 14458 57468 14464 57520
rect 14516 57508 14522 57520
rect 75546 57508 75552 57520
rect 14516 57480 75552 57508
rect 14516 57468 14522 57480
rect 75546 57468 75552 57480
rect 75604 57468 75610 57520
rect 75822 57468 75828 57520
rect 75880 57508 75886 57520
rect 148686 57508 148692 57520
rect 75880 57480 148692 57508
rect 75880 57468 75886 57480
rect 148686 57468 148692 57480
rect 148744 57468 148750 57520
rect 162118 57468 162124 57520
rect 162176 57508 162182 57520
rect 171318 57508 171324 57520
rect 162176 57480 171324 57508
rect 162176 57468 162182 57480
rect 171318 57468 171324 57480
rect 171376 57468 171382 57520
rect 183002 57468 183008 57520
rect 183060 57508 183066 57520
rect 184198 57508 184204 57520
rect 183060 57480 184204 57508
rect 183060 57468 183066 57480
rect 184198 57468 184204 57480
rect 184256 57468 184262 57520
rect 235442 57468 235448 57520
rect 235500 57508 235506 57520
rect 384301 57511 384359 57517
rect 384301 57508 384313 57511
rect 235500 57480 384313 57508
rect 235500 57468 235506 57480
rect 384301 57477 384313 57480
rect 384347 57477 384359 57511
rect 384301 57471 384359 57477
rect 384390 57468 384396 57520
rect 384448 57508 384454 57520
rect 384942 57508 384948 57520
rect 384448 57480 384948 57508
rect 384448 57468 384454 57480
rect 384942 57468 384948 57480
rect 385000 57468 385006 57520
rect 385310 57468 385316 57520
rect 385368 57508 385374 57520
rect 386322 57508 386328 57520
rect 385368 57480 386328 57508
rect 385368 57468 385374 57480
rect 386322 57468 386328 57480
rect 386380 57468 386386 57520
rect 387150 57468 387156 57520
rect 387208 57508 387214 57520
rect 387702 57508 387708 57520
rect 387208 57480 387708 57508
rect 387208 57468 387214 57480
rect 387702 57468 387708 57480
rect 387760 57468 387766 57520
rect 387978 57468 387984 57520
rect 388036 57508 388042 57520
rect 389082 57508 389088 57520
rect 388036 57480 389088 57508
rect 388036 57468 388042 57480
rect 389082 57468 389088 57480
rect 389140 57468 389146 57520
rect 389818 57468 389824 57520
rect 389876 57508 389882 57520
rect 390462 57508 390468 57520
rect 389876 57480 390468 57508
rect 389876 57468 389882 57480
rect 390462 57468 390468 57480
rect 390520 57468 390526 57520
rect 390738 57468 390744 57520
rect 390796 57508 390802 57520
rect 391842 57508 391848 57520
rect 390796 57480 391848 57508
rect 390796 57468 390802 57480
rect 391842 57468 391848 57480
rect 391900 57468 391906 57520
rect 392578 57468 392584 57520
rect 392636 57508 392642 57520
rect 393222 57508 393228 57520
rect 392636 57480 393228 57508
rect 392636 57468 392642 57480
rect 393222 57468 393228 57480
rect 393280 57468 393286 57520
rect 393406 57468 393412 57520
rect 393464 57508 393470 57520
rect 394602 57508 394608 57520
rect 393464 57480 394608 57508
rect 393464 57468 393470 57480
rect 394602 57468 394608 57480
rect 394660 57468 394666 57520
rect 395246 57468 395252 57520
rect 395304 57508 395310 57520
rect 395982 57508 395988 57520
rect 395304 57480 395988 57508
rect 395304 57468 395310 57480
rect 395982 57468 395988 57480
rect 396040 57468 396046 57520
rect 396166 57468 396172 57520
rect 396224 57508 396230 57520
rect 397270 57508 397276 57520
rect 396224 57480 397276 57508
rect 396224 57468 396230 57480
rect 397270 57468 397276 57480
rect 397328 57468 397334 57520
rect 398006 57468 398012 57520
rect 398064 57508 398070 57520
rect 398742 57508 398748 57520
rect 398064 57480 398748 57508
rect 398064 57468 398070 57480
rect 398742 57468 398748 57480
rect 398800 57468 398806 57520
rect 400858 57468 400864 57520
rect 400916 57508 400922 57520
rect 401594 57508 401600 57520
rect 400916 57480 401600 57508
rect 400916 57468 400922 57480
rect 401594 57468 401600 57480
rect 401652 57468 401658 57520
rect 401686 57468 401692 57520
rect 401744 57508 401750 57520
rect 464617 57511 464675 57517
rect 464617 57508 464629 57511
rect 401744 57480 464629 57508
rect 401744 57468 401750 57480
rect 464617 57477 464629 57480
rect 464663 57477 464675 57511
rect 464617 57471 464675 57477
rect 466546 57468 466552 57520
rect 466604 57508 466610 57520
rect 467466 57508 467472 57520
rect 466604 57480 467472 57508
rect 466604 57468 466610 57480
rect 467466 57468 467472 57480
rect 467524 57468 467530 57520
rect 469122 57468 469128 57520
rect 469180 57508 469186 57520
rect 485498 57508 485504 57520
rect 469180 57480 485504 57508
rect 469180 57468 469186 57480
rect 485498 57468 485504 57480
rect 485556 57468 485562 57520
rect 18598 57400 18604 57452
rect 18656 57440 18662 57452
rect 134242 57440 134248 57452
rect 18656 57412 134248 57440
rect 18656 57400 18662 57412
rect 134242 57400 134248 57412
rect 134300 57400 134306 57452
rect 161382 57400 161388 57452
rect 161440 57440 161446 57452
rect 176654 57440 176660 57452
rect 161440 57412 176660 57440
rect 161440 57400 161446 57412
rect 176654 57400 176660 57412
rect 176712 57400 176718 57452
rect 177298 57400 177304 57452
rect 177356 57440 177362 57452
rect 179414 57440 179420 57452
rect 177356 57412 179420 57440
rect 177356 57400 177362 57412
rect 179414 57400 179420 57412
rect 179472 57400 179478 57452
rect 219158 57400 219164 57452
rect 219216 57440 219222 57452
rect 222838 57440 222844 57452
rect 219216 57412 222844 57440
rect 219216 57400 219222 57412
rect 222838 57400 222844 57412
rect 222896 57400 222902 57452
rect 238110 57400 238116 57452
rect 238168 57440 238174 57452
rect 238662 57440 238668 57452
rect 238168 57412 238668 57440
rect 238168 57400 238174 57412
rect 238662 57400 238668 57412
rect 238720 57400 238726 57452
rect 240870 57400 240876 57452
rect 240928 57440 240934 57452
rect 241422 57440 241428 57452
rect 240928 57412 241428 57440
rect 240928 57400 240934 57412
rect 241422 57400 241428 57412
rect 241480 57400 241486 57452
rect 241698 57400 241704 57452
rect 241756 57440 241762 57452
rect 242802 57440 242808 57452
rect 241756 57412 242808 57440
rect 241756 57400 241762 57412
rect 242802 57400 242808 57412
rect 242860 57400 242866 57452
rect 243538 57400 243544 57452
rect 243596 57440 243602 57452
rect 244182 57440 244188 57452
rect 243596 57412 244188 57440
rect 243596 57400 243602 57412
rect 244182 57400 244188 57412
rect 244240 57400 244246 57452
rect 244458 57400 244464 57452
rect 244516 57440 244522 57452
rect 245470 57440 245476 57452
rect 244516 57412 245476 57440
rect 244516 57400 244522 57412
rect 245470 57400 245476 57412
rect 245528 57400 245534 57452
rect 246206 57400 246212 57452
rect 246264 57440 246270 57452
rect 246942 57440 246948 57452
rect 246264 57412 246948 57440
rect 246264 57400 246270 57412
rect 246942 57400 246948 57412
rect 247000 57400 247006 57452
rect 407758 57440 407764 57452
rect 247052 57412 407764 57440
rect 29638 57332 29644 57384
rect 29696 57372 29702 57384
rect 164970 57372 164976 57384
rect 29696 57344 164976 57372
rect 29696 57332 29702 57344
rect 164970 57332 164976 57344
rect 165028 57332 165034 57384
rect 188430 57332 188436 57384
rect 188488 57372 188494 57384
rect 196618 57372 196624 57384
rect 188488 57344 196624 57372
rect 188488 57332 188494 57344
rect 196618 57332 196624 57344
rect 196676 57332 196682 57384
rect 233602 57332 233608 57384
rect 233660 57372 233666 57384
rect 238205 57375 238263 57381
rect 238205 57372 238217 57375
rect 233660 57344 238217 57372
rect 233660 57332 233666 57344
rect 238205 57341 238217 57344
rect 238251 57341 238263 57375
rect 238205 57335 238263 57341
rect 239950 57332 239956 57384
rect 240008 57372 240014 57384
rect 247052 57372 247080 57412
rect 407758 57400 407764 57412
rect 407816 57400 407822 57452
rect 410518 57400 410524 57452
rect 410576 57440 410582 57452
rect 423214 57440 423220 57452
rect 410576 57412 423220 57440
rect 410576 57400 410582 57412
rect 423214 57400 423220 57412
rect 423272 57400 423278 57452
rect 423582 57400 423588 57452
rect 423640 57440 423646 57452
rect 473814 57440 473820 57452
rect 423640 57412 473820 57440
rect 423640 57400 423646 57412
rect 473814 57400 473820 57412
rect 473872 57400 473878 57452
rect 476022 57400 476028 57452
rect 476080 57440 476086 57452
rect 487338 57440 487344 57452
rect 476080 57412 487344 57440
rect 476080 57400 476086 57412
rect 487338 57400 487344 57412
rect 487396 57400 487402 57452
rect 512638 57400 512644 57452
rect 512696 57440 512702 57452
rect 513282 57440 513288 57452
rect 512696 57412 513288 57440
rect 512696 57400 512702 57412
rect 513282 57400 513288 57412
rect 513340 57400 513346 57452
rect 240008 57344 247080 57372
rect 240008 57332 240014 57344
rect 247126 57332 247132 57384
rect 247184 57372 247190 57384
rect 248322 57372 248328 57384
rect 247184 57344 248328 57372
rect 247184 57332 247190 57344
rect 248322 57332 248328 57344
rect 248380 57332 248386 57384
rect 248966 57332 248972 57384
rect 249024 57372 249030 57384
rect 249702 57372 249708 57384
rect 249024 57344 249708 57372
rect 249024 57332 249030 57344
rect 249702 57332 249708 57344
rect 249760 57332 249766 57384
rect 249886 57332 249892 57384
rect 249944 57372 249950 57384
rect 250990 57372 250996 57384
rect 249944 57344 250996 57372
rect 249944 57332 249950 57344
rect 250990 57332 250996 57344
rect 251048 57332 251054 57384
rect 251634 57332 251640 57384
rect 251692 57372 251698 57384
rect 252462 57372 252468 57384
rect 251692 57344 252468 57372
rect 251692 57332 251698 57344
rect 252462 57332 252468 57344
rect 252520 57332 252526 57384
rect 252554 57332 252560 57384
rect 252612 57372 252618 57384
rect 253750 57372 253756 57384
rect 252612 57344 253756 57372
rect 252612 57332 252618 57344
rect 253750 57332 253756 57344
rect 253808 57332 253814 57384
rect 254394 57332 254400 57384
rect 254452 57372 254458 57384
rect 255222 57372 255228 57384
rect 254452 57344 255228 57372
rect 254452 57332 254458 57344
rect 255222 57332 255228 57344
rect 255280 57332 255286 57384
rect 255314 57332 255320 57384
rect 255372 57372 255378 57384
rect 256602 57372 256608 57384
rect 255372 57344 256608 57372
rect 255372 57332 255378 57344
rect 256602 57332 256608 57344
rect 256660 57332 256666 57384
rect 257982 57332 257988 57384
rect 258040 57372 258046 57384
rect 446033 57375 446091 57381
rect 446033 57372 446045 57375
rect 258040 57344 446045 57372
rect 258040 57332 258046 57344
rect 446033 57341 446045 57344
rect 446079 57341 446091 57375
rect 446033 57335 446091 57341
rect 448422 57332 448428 57384
rect 448480 57372 448486 57384
rect 449437 57375 449495 57381
rect 449437 57372 449449 57375
rect 448480 57344 449449 57372
rect 448480 57332 448486 57344
rect 449437 57341 449449 57344
rect 449483 57341 449495 57375
rect 449437 57335 449495 57341
rect 455322 57332 455328 57384
rect 455380 57372 455386 57384
rect 481910 57372 481916 57384
rect 455380 57344 481916 57372
rect 455380 57332 455386 57344
rect 481910 57332 481916 57344
rect 481968 57332 481974 57384
rect 22738 57264 22744 57316
rect 22796 57304 22802 57316
rect 163130 57304 163136 57316
rect 22796 57276 163136 57304
rect 22796 57264 22802 57276
rect 163130 57264 163136 57276
rect 163188 57264 163194 57316
rect 165522 57264 165528 57316
rect 165580 57304 165586 57316
rect 177574 57304 177580 57316
rect 165580 57276 177580 57304
rect 165580 57264 165586 57276
rect 177574 57264 177580 57276
rect 177632 57264 177638 57316
rect 190270 57264 190276 57316
rect 190328 57304 190334 57316
rect 202138 57304 202144 57316
rect 190328 57276 202144 57304
rect 190328 57264 190334 57276
rect 202138 57264 202144 57276
rect 202196 57264 202202 57316
rect 208210 57264 208216 57316
rect 208268 57304 208274 57316
rect 258718 57304 258724 57316
rect 208268 57276 258724 57304
rect 208268 57264 208274 57276
rect 258718 57264 258724 57276
rect 258776 57264 258782 57316
rect 258902 57264 258908 57316
rect 258960 57304 258966 57316
rect 259362 57304 259368 57316
rect 258960 57276 259368 57304
rect 258960 57264 258966 57276
rect 259362 57264 259368 57276
rect 259420 57264 259426 57316
rect 261570 57264 261576 57316
rect 261628 57304 261634 57316
rect 489178 57304 489184 57316
rect 261628 57276 264376 57304
rect 261628 57264 261634 57276
rect 7558 57196 7564 57248
rect 7616 57236 7622 57248
rect 166718 57236 166724 57248
rect 7616 57208 166724 57236
rect 7616 57196 7622 57208
rect 166718 57196 166724 57208
rect 166776 57196 166782 57248
rect 183922 57196 183928 57248
rect 183980 57236 183986 57248
rect 188430 57236 188436 57248
rect 183980 57208 188436 57236
rect 183980 57196 183986 57208
rect 188430 57196 188436 57208
rect 188488 57196 188494 57248
rect 189350 57196 189356 57248
rect 189408 57236 189414 57248
rect 204898 57236 204904 57248
rect 189408 57208 204904 57236
rect 189408 57196 189414 57208
rect 204898 57196 204904 57208
rect 204956 57196 204962 57248
rect 210142 57196 210148 57248
rect 210200 57236 210206 57248
rect 264238 57236 264244 57248
rect 210200 57208 264244 57236
rect 210200 57196 210206 57208
rect 264238 57196 264244 57208
rect 264296 57196 264302 57248
rect 264348 57236 264376 57276
rect 264992 57276 489184 57304
rect 264992 57236 265020 57276
rect 489178 57264 489184 57276
rect 489236 57264 489242 57316
rect 264348 57208 265020 57236
rect 265250 57196 265256 57248
rect 265308 57236 265314 57248
rect 507118 57236 507124 57248
rect 265308 57208 507124 57236
rect 265308 57196 265314 57208
rect 507118 57196 507124 57208
rect 507176 57196 507182 57248
rect 68278 57128 68284 57180
rect 68336 57168 68342 57180
rect 84562 57168 84568 57180
rect 68336 57140 84568 57168
rect 68336 57128 68342 57140
rect 84562 57128 84568 57140
rect 84620 57128 84626 57180
rect 211982 57128 211988 57180
rect 212040 57168 212046 57180
rect 275281 57171 275339 57177
rect 275281 57168 275293 57171
rect 212040 57140 275293 57168
rect 212040 57128 212046 57140
rect 275281 57137 275293 57140
rect 275327 57137 275339 57171
rect 275281 57131 275339 57137
rect 275388 57140 282914 57168
rect 69658 57060 69664 57112
rect 69716 57100 69722 57112
rect 83642 57100 83648 57112
rect 69716 57072 83648 57100
rect 69716 57060 69722 57072
rect 83642 57060 83648 57072
rect 83700 57060 83706 57112
rect 257062 57060 257068 57112
rect 257120 57100 257126 57112
rect 257982 57100 257988 57112
rect 257120 57072 257988 57100
rect 257120 57060 257126 57072
rect 257982 57060 257988 57072
rect 258040 57060 258046 57112
rect 262858 57060 262864 57112
rect 262916 57100 262922 57112
rect 275388 57100 275416 57140
rect 262916 57072 275416 57100
rect 282886 57100 282914 57140
rect 287698 57128 287704 57180
rect 287756 57168 287762 57180
rect 293218 57168 293224 57180
rect 287756 57140 293224 57168
rect 287756 57128 287762 57140
rect 293218 57128 293224 57140
rect 293276 57128 293282 57180
rect 342898 57128 342904 57180
rect 342956 57168 342962 57180
rect 344005 57171 344063 57177
rect 344005 57168 344017 57171
rect 342956 57140 344017 57168
rect 342956 57128 342962 57140
rect 344005 57137 344017 57140
rect 344051 57137 344063 57171
rect 344005 57131 344063 57137
rect 364429 57171 364487 57177
rect 364429 57137 364441 57171
rect 364475 57168 364487 57171
rect 371878 57168 371884 57180
rect 364475 57140 371884 57168
rect 364475 57137 364487 57140
rect 364429 57131 364487 57137
rect 371878 57128 371884 57140
rect 371936 57128 371942 57180
rect 384301 57171 384359 57177
rect 384301 57137 384313 57171
rect 384347 57168 384359 57171
rect 389818 57168 389824 57180
rect 384347 57140 389824 57168
rect 384347 57137 384359 57140
rect 384301 57131 384359 57137
rect 389818 57128 389824 57140
rect 389876 57128 389882 57180
rect 446033 57171 446091 57177
rect 446033 57137 446045 57171
rect 446079 57168 446091 57171
rect 450538 57168 450544 57180
rect 446079 57140 450544 57168
rect 446079 57137 446091 57140
rect 446033 57131 446091 57137
rect 450538 57128 450544 57140
rect 450596 57128 450602 57180
rect 462222 57128 462228 57180
rect 462280 57168 462286 57180
rect 468481 57171 468539 57177
rect 468481 57168 468493 57171
rect 462280 57140 468493 57168
rect 462280 57128 462286 57140
rect 468481 57137 468493 57140
rect 468527 57137 468539 57171
rect 468481 57131 468539 57137
rect 473262 57128 473268 57180
rect 473320 57168 473326 57180
rect 486418 57168 486424 57180
rect 473320 57140 486424 57168
rect 473320 57128 473326 57140
rect 486418 57128 486424 57140
rect 486476 57128 486482 57180
rect 504542 57128 504548 57180
rect 504600 57168 504606 57180
rect 505002 57168 505008 57180
rect 504600 57140 505008 57168
rect 504600 57128 504606 57140
rect 505002 57128 505008 57140
rect 505060 57128 505066 57180
rect 315758 57100 315764 57112
rect 282886 57072 315764 57100
rect 262916 57060 262922 57072
rect 315758 57060 315764 57072
rect 315816 57060 315822 57112
rect 471793 57103 471851 57109
rect 471793 57069 471805 57103
rect 471839 57100 471851 57103
rect 480070 57100 480076 57112
rect 471839 57072 480076 57100
rect 471839 57069 471851 57072
rect 471793 57063 471851 57069
rect 480070 57060 480076 57072
rect 480128 57060 480134 57112
rect 71774 56992 71780 57044
rect 71832 57032 71838 57044
rect 81894 57032 81900 57044
rect 71832 57004 81900 57032
rect 71832 56992 71838 57004
rect 81894 56992 81900 57004
rect 81952 56992 81958 57044
rect 239030 56992 239036 57044
rect 239088 57032 239094 57044
rect 246298 57032 246304 57044
rect 239088 57004 246304 57032
rect 239088 56992 239094 57004
rect 246298 56992 246304 57004
rect 246356 56992 246362 57044
rect 264330 56992 264336 57044
rect 264388 57032 264394 57044
rect 264882 57032 264888 57044
rect 264388 57004 264888 57032
rect 264388 56992 264394 57004
rect 264882 56992 264888 57004
rect 264940 56992 264946 57044
rect 266998 56992 267004 57044
rect 267056 57032 267062 57044
rect 267642 57032 267648 57044
rect 267056 57004 267648 57032
rect 267056 56992 267062 57004
rect 267642 56992 267648 57004
rect 267700 56992 267706 57044
rect 267918 56992 267924 57044
rect 267976 57032 267982 57044
rect 269022 57032 269028 57044
rect 267976 57004 269028 57032
rect 267976 56992 267982 57004
rect 269022 56992 269028 57004
rect 269080 56992 269086 57044
rect 269758 56992 269764 57044
rect 269816 57032 269822 57044
rect 270402 57032 270408 57044
rect 269816 57004 270408 57032
rect 269816 56992 269822 57004
rect 270402 56992 270408 57004
rect 270460 56992 270466 57044
rect 270678 56992 270684 57044
rect 270736 57032 270742 57044
rect 271690 57032 271696 57044
rect 270736 57004 271696 57032
rect 270736 56992 270742 57004
rect 271690 56992 271696 57004
rect 271748 56992 271754 57044
rect 272426 56992 272432 57044
rect 272484 57032 272490 57044
rect 273162 57032 273168 57044
rect 272484 57004 273168 57032
rect 272484 56992 272490 57004
rect 273162 56992 273168 57004
rect 273220 56992 273226 57044
rect 320174 57032 320180 57044
rect 287026 57004 320180 57032
rect 65610 56924 65616 56976
rect 65668 56964 65674 56976
rect 72513 56967 72571 56973
rect 72513 56964 72525 56967
rect 65668 56936 72525 56964
rect 65668 56924 65674 56936
rect 72513 56933 72525 56936
rect 72559 56933 72571 56967
rect 72513 56927 72571 56933
rect 278130 56924 278136 56976
rect 278188 56964 278194 56976
rect 287026 56964 287054 57004
rect 320174 56992 320180 57004
rect 320232 56992 320238 57044
rect 502702 56992 502708 57044
rect 502760 57032 502766 57044
rect 503530 57032 503536 57044
rect 502760 57004 503536 57032
rect 502760 56992 502766 57004
rect 503530 56992 503536 57004
rect 503588 56992 503594 57044
rect 278188 56936 287054 56964
rect 278188 56924 278194 56936
rect 275281 56899 275339 56905
rect 275281 56865 275293 56899
rect 275327 56896 275339 56899
rect 284938 56896 284944 56908
rect 275327 56868 284944 56896
rect 275327 56865 275339 56868
rect 275281 56859 275339 56865
rect 284938 56856 284944 56868
rect 284996 56856 285002 56908
rect 316678 56856 316684 56908
rect 316736 56896 316742 56908
rect 319346 56896 319352 56908
rect 316736 56868 319352 56896
rect 316736 56856 316742 56868
rect 319346 56856 319352 56868
rect 319404 56856 319410 56908
rect 86218 56788 86224 56840
rect 86276 56828 86282 56840
rect 89990 56828 89996 56840
rect 86276 56800 89996 56828
rect 86276 56788 86282 56800
rect 89990 56788 89996 56800
rect 90048 56788 90054 56840
rect 186682 56720 186688 56772
rect 186740 56760 186746 56772
rect 191098 56760 191104 56772
rect 186740 56732 191104 56760
rect 186740 56720 186746 56732
rect 191098 56720 191104 56732
rect 191156 56720 191162 56772
rect 220998 56720 221004 56772
rect 221056 56760 221062 56772
rect 228358 56760 228364 56772
rect 221056 56732 228364 56760
rect 221056 56720 221062 56732
rect 228358 56720 228364 56732
rect 228416 56720 228422 56772
rect 237190 56652 237196 56704
rect 237248 56692 237254 56704
rect 240778 56692 240784 56704
rect 237248 56664 240784 56692
rect 237248 56652 237254 56664
rect 240778 56652 240784 56664
rect 240836 56652 240842 56704
rect 373626 56652 373632 56704
rect 373684 56692 373690 56704
rect 374638 56692 374644 56704
rect 373684 56664 374644 56692
rect 373684 56652 373690 56664
rect 374638 56652 374644 56664
rect 374696 56652 374702 56704
rect 102686 56584 102692 56636
rect 102744 56624 102750 56636
rect 105538 56624 105544 56636
rect 102744 56596 105544 56624
rect 102744 56584 102750 56596
rect 105538 56584 105544 56596
rect 105596 56584 105602 56636
rect 170398 56584 170404 56636
rect 170456 56624 170462 56636
rect 172146 56624 172152 56636
rect 170456 56596 172152 56624
rect 170456 56584 170462 56596
rect 172146 56584 172152 56596
rect 172204 56584 172210 56636
rect 179322 56584 179328 56636
rect 179380 56624 179386 56636
rect 181254 56624 181260 56636
rect 179380 56596 181260 56624
rect 179380 56584 179386 56596
rect 181254 56584 181260 56596
rect 181312 56584 181318 56636
rect 218238 56584 218244 56636
rect 218296 56624 218302 56636
rect 220078 56624 220084 56636
rect 218296 56596 220084 56624
rect 218296 56584 218302 56596
rect 220078 56584 220084 56596
rect 220136 56584 220142 56636
rect 273346 56584 273352 56636
rect 273404 56624 273410 56636
rect 274450 56624 274456 56636
rect 273404 56596 274456 56624
rect 273404 56584 273410 56596
rect 274450 56584 274456 56596
rect 274508 56584 274514 56636
rect 275186 56584 275192 56636
rect 275244 56624 275250 56636
rect 275922 56624 275928 56636
rect 275244 56596 275928 56624
rect 275244 56584 275250 56596
rect 275922 56584 275928 56596
rect 275980 56584 275986 56636
rect 276014 56584 276020 56636
rect 276072 56624 276078 56636
rect 277302 56624 277308 56636
rect 276072 56596 277308 56624
rect 276072 56584 276078 56596
rect 277302 56584 277308 56596
rect 277360 56584 277366 56636
rect 277854 56584 277860 56636
rect 277912 56624 277918 56636
rect 278682 56624 278688 56636
rect 277912 56596 278688 56624
rect 277912 56584 277918 56596
rect 278682 56584 278688 56596
rect 278740 56584 278746 56636
rect 278774 56584 278780 56636
rect 278832 56624 278838 56636
rect 280062 56624 280068 56636
rect 278832 56596 280068 56624
rect 278832 56584 278838 56596
rect 280062 56584 280068 56596
rect 280120 56584 280126 56636
rect 280522 56584 280528 56636
rect 280580 56624 280586 56636
rect 281350 56624 281356 56636
rect 280580 56596 281356 56624
rect 280580 56584 280586 56596
rect 281350 56584 281356 56596
rect 281408 56584 281414 56636
rect 282362 56584 282368 56636
rect 282420 56624 282426 56636
rect 282822 56624 282828 56636
rect 282420 56596 282828 56624
rect 282420 56584 282426 56596
rect 282822 56584 282828 56596
rect 282880 56584 282886 56636
rect 295978 56584 295984 56636
rect 296036 56624 296042 56636
rect 296806 56624 296812 56636
rect 296036 56596 296812 56624
rect 296036 56584 296042 56596
rect 296806 56584 296812 56596
rect 296864 56584 296870 56636
rect 421558 56584 421564 56636
rect 421616 56624 421622 56636
rect 422294 56624 422300 56636
rect 421616 56596 422300 56624
rect 421616 56584 421622 56596
rect 422294 56584 422300 56596
rect 422352 56584 422358 56636
rect 487062 56584 487068 56636
rect 487120 56624 487126 56636
rect 490006 56624 490012 56636
rect 487120 56596 490012 56624
rect 487120 56584 487126 56596
rect 490006 56584 490012 56596
rect 490064 56584 490070 56636
rect 62022 56380 62028 56432
rect 62080 56420 62086 56432
rect 87322 56420 87328 56432
rect 62080 56392 87328 56420
rect 62080 56380 62086 56392
rect 87322 56380 87328 56392
rect 87380 56380 87386 56432
rect 41322 56312 41328 56364
rect 41380 56352 41386 56364
rect 71774 56352 71780 56364
rect 41380 56324 71780 56352
rect 41380 56312 41386 56324
rect 71774 56312 71780 56324
rect 71832 56312 71838 56364
rect 37182 56244 37188 56296
rect 37240 56284 37246 56296
rect 80974 56284 80980 56296
rect 37240 56256 80980 56284
rect 37240 56244 37246 56256
rect 80974 56244 80980 56256
rect 81032 56244 81038 56296
rect 345658 56244 345664 56296
rect 345716 56284 345722 56296
rect 452102 56284 452108 56296
rect 345716 56256 452108 56284
rect 345716 56244 345722 56256
rect 452102 56244 452108 56256
rect 452160 56244 452166 56296
rect 34422 56176 34428 56228
rect 34480 56216 34486 56228
rect 79962 56216 79968 56228
rect 34480 56188 79968 56216
rect 34480 56176 34486 56188
rect 79962 56176 79968 56188
rect 80020 56176 80026 56228
rect 188338 56176 188344 56228
rect 188396 56216 188402 56228
rect 297726 56216 297732 56228
rect 188396 56188 297732 56216
rect 188396 56176 188402 56188
rect 297726 56176 297732 56188
rect 297784 56176 297790 56228
rect 380802 56176 380808 56228
rect 380860 56216 380866 56228
rect 501598 56216 501604 56228
rect 380860 56188 501604 56216
rect 380860 56176 380866 56188
rect 501598 56176 501604 56188
rect 501656 56176 501662 56228
rect 22002 56108 22008 56160
rect 22060 56148 22066 56160
rect 77202 56148 77208 56160
rect 22060 56120 77208 56148
rect 22060 56108 22066 56120
rect 77202 56108 77208 56120
rect 77260 56108 77266 56160
rect 282178 56108 282184 56160
rect 282236 56148 282242 56160
rect 434070 56148 434076 56160
rect 282236 56120 434076 56148
rect 282236 56108 282242 56120
rect 434070 56108 434076 56120
rect 434128 56108 434134 56160
rect 43438 56040 43444 56092
rect 43496 56080 43502 56092
rect 109034 56080 109040 56092
rect 43496 56052 109040 56080
rect 43496 56040 43502 56052
rect 109034 56040 109040 56052
rect 109092 56040 109098 56092
rect 260098 56040 260104 56092
rect 260156 56080 260162 56092
rect 427722 56080 427728 56092
rect 260156 56052 427728 56080
rect 260156 56040 260162 56052
rect 427722 56040 427728 56052
rect 427780 56040 427786 56092
rect 25498 55972 25504 56024
rect 25556 56012 25562 56024
rect 103514 56012 103520 56024
rect 25556 55984 103520 56012
rect 25556 55972 25562 55984
rect 103514 55972 103520 55984
rect 103572 55972 103578 56024
rect 249058 55972 249064 56024
rect 249116 56012 249122 56024
rect 426802 56012 426808 56024
rect 249116 55984 426808 56012
rect 249116 55972 249122 55984
rect 426802 55972 426808 55984
rect 426860 55972 426866 56024
rect 65518 55904 65524 55956
rect 65576 55944 65582 55956
rect 146018 55944 146024 55956
rect 65576 55916 146024 55944
rect 65576 55904 65582 55916
rect 146018 55904 146024 55916
rect 146076 55904 146082 55956
rect 262490 55904 262496 55956
rect 262548 55944 262554 55956
rect 483658 55944 483664 55956
rect 262548 55916 483664 55944
rect 262548 55904 262554 55916
rect 483658 55904 483664 55916
rect 483716 55904 483722 55956
rect 58618 55836 58624 55888
rect 58676 55876 58682 55888
rect 142338 55876 142344 55888
rect 58676 55848 142344 55876
rect 58676 55836 58682 55848
rect 142338 55836 142344 55848
rect 142396 55836 142402 55888
rect 259822 55836 259828 55888
rect 259880 55876 259886 55888
rect 485038 55876 485044 55888
rect 259880 55848 485044 55876
rect 259880 55836 259886 55848
rect 485038 55836 485044 55848
rect 485096 55836 485102 55888
rect 47578 54680 47584 54732
rect 47636 54720 47642 54732
rect 110506 54720 110512 54732
rect 47636 54692 110512 54720
rect 47636 54680 47642 54692
rect 110506 54680 110512 54692
rect 110564 54680 110570 54732
rect 39298 54612 39304 54664
rect 39356 54652 39362 54664
rect 106366 54652 106372 54664
rect 39356 54624 106372 54652
rect 39356 54612 39362 54624
rect 106366 54612 106372 54624
rect 106424 54612 106430 54664
rect 35158 54544 35164 54596
rect 35216 54584 35222 54596
rect 104894 54584 104900 54596
rect 35216 54556 104900 54584
rect 35216 54544 35222 54556
rect 104894 54544 104900 54556
rect 104952 54544 104958 54596
rect 318058 54544 318064 54596
rect 318116 54584 318122 54596
rect 440510 54584 440516 54596
rect 318116 54556 440516 54584
rect 318116 54544 318122 54556
rect 440510 54544 440516 54556
rect 440568 54544 440574 54596
rect 15838 54476 15844 54528
rect 15896 54516 15902 54528
rect 132586 54516 132592 54528
rect 15896 54488 132592 54516
rect 15896 54476 15902 54488
rect 132586 54476 132592 54488
rect 132644 54476 132650 54528
rect 251818 54476 251824 54528
rect 251876 54516 251882 54528
rect 429286 54516 429292 54528
rect 251876 54488 429292 54516
rect 251876 54476 251882 54488
rect 429286 54476 429292 54488
rect 429344 54476 429350 54528
rect 519814 46860 519820 46912
rect 519872 46900 519878 46912
rect 580166 46900 580172 46912
rect 519872 46872 580172 46900
rect 519872 46860 519878 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 266998 37884 267004 37936
rect 267056 37924 267062 37936
rect 429194 37924 429200 37936
rect 267056 37896 429200 37924
rect 267056 37884 267062 37896
rect 429194 37884 429200 37896
rect 429252 37884 429258 37936
rect 142062 36524 142068 36576
rect 142120 36564 142126 36576
rect 285766 36564 285772 36576
rect 142120 36536 285772 36564
rect 142120 36524 142126 36536
rect 285766 36524 285772 36536
rect 285824 36524 285830 36576
rect 286318 36524 286324 36576
rect 286376 36564 286382 36576
rect 432046 36564 432052 36576
rect 286376 36536 432052 36564
rect 286376 36524 286382 36536
rect 432046 36524 432052 36536
rect 432104 36524 432110 36576
rect 233878 33736 233884 33788
rect 233936 33776 233942 33788
rect 425146 33776 425152 33788
rect 233936 33748 425152 33776
rect 233936 33736 233942 33748
rect 425146 33736 425152 33748
rect 425204 33736 425210 33788
rect 519722 33056 519728 33108
rect 519780 33096 519786 33108
rect 580166 33096 580172 33108
rect 519780 33068 580172 33096
rect 519780 33056 519786 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 160002 32376 160008 32428
rect 160060 32416 160066 32428
rect 291286 32416 291292 32428
rect 160060 32388 291292 32416
rect 160060 32376 160066 32388
rect 291286 32376 291292 32388
rect 291344 32376 291350 32428
rect 360838 32376 360844 32428
rect 360896 32416 360902 32428
rect 449894 32416 449900 32428
rect 360896 32388 449900 32416
rect 360896 32376 360902 32388
rect 449894 32376 449900 32388
rect 449952 32376 449958 32428
rect 153102 31016 153108 31068
rect 153160 31056 153166 31068
rect 288526 31056 288532 31068
rect 153160 31028 288532 31056
rect 153160 31016 153166 31028
rect 288526 31016 288532 31028
rect 288584 31016 288590 31068
rect 320818 31016 320824 31068
rect 320876 31056 320882 31068
rect 443086 31056 443092 31068
rect 320876 31028 443092 31056
rect 320876 31016 320882 31028
rect 443086 31016 443092 31028
rect 443144 31016 443150 31068
rect 61930 29588 61936 29640
rect 61988 29628 61994 29640
rect 144178 29628 144184 29640
rect 61988 29600 144184 29628
rect 61988 29588 61994 29600
rect 144178 29588 144184 29600
rect 144236 29588 144242 29640
rect 209038 29588 209044 29640
rect 209096 29628 209102 29640
rect 299566 29628 299572 29640
rect 209096 29600 299572 29628
rect 209096 29588 209102 29600
rect 299566 29588 299572 29600
rect 299624 29588 299630 29640
rect 374638 29588 374644 29640
rect 374696 29628 374702 29640
rect 481634 29628 481640 29640
rect 374696 29600 481640 29628
rect 374696 29588 374702 29600
rect 481634 29588 481640 29600
rect 481692 29588 481698 29640
rect 144822 28228 144828 28280
rect 144880 28268 144886 28280
rect 170398 28268 170404 28280
rect 144880 28240 170404 28268
rect 144880 28228 144886 28240
rect 170398 28228 170404 28240
rect 170456 28228 170462 28280
rect 289170 28228 289176 28280
rect 289228 28268 289234 28280
rect 434806 28268 434812 28280
rect 289228 28240 434812 28268
rect 289228 28228 289234 28240
rect 434806 28228 434812 28240
rect 434864 28228 434870 28280
rect 173802 26868 173808 26920
rect 173860 26908 173866 26920
rect 294046 26908 294052 26920
rect 173860 26880 294052 26908
rect 173860 26868 173866 26880
rect 294046 26868 294052 26880
rect 294104 26868 294110 26920
rect 300118 26868 300124 26920
rect 300176 26908 300182 26920
rect 441614 26908 441620 26920
rect 300176 26880 441620 26908
rect 300176 26868 300182 26880
rect 441614 26868 441620 26880
rect 441672 26868 441678 26920
rect 51718 25508 51724 25560
rect 51776 25548 51782 25560
rect 111794 25548 111800 25560
rect 51776 25520 111800 25548
rect 51776 25508 51782 25520
rect 111794 25508 111800 25520
rect 111852 25508 111858 25560
rect 113082 25508 113088 25560
rect 113140 25548 113146 25560
rect 129826 25548 129832 25560
rect 113140 25520 129832 25548
rect 113140 25508 113146 25520
rect 129826 25508 129832 25520
rect 129884 25508 129890 25560
rect 222838 25508 222844 25560
rect 222896 25548 222902 25560
rect 327166 25548 327172 25560
rect 222896 25520 327172 25548
rect 222896 25508 222902 25520
rect 327166 25508 327172 25520
rect 327224 25508 327230 25560
rect 376570 25508 376576 25560
rect 376628 25548 376634 25560
rect 486418 25548 486424 25560
rect 376628 25520 486424 25548
rect 376628 25508 376634 25520
rect 486418 25508 486424 25520
rect 486476 25508 486482 25560
rect 81342 24080 81348 24132
rect 81400 24120 81406 24132
rect 121454 24120 121460 24132
rect 81400 24092 121460 24120
rect 81400 24080 81406 24092
rect 121454 24080 121460 24092
rect 121512 24080 121518 24132
rect 241422 24080 241428 24132
rect 241480 24120 241486 24132
rect 412726 24120 412732 24132
rect 241480 24092 412732 24120
rect 241480 24080 241486 24092
rect 412726 24080 412732 24092
rect 412784 24080 412790 24132
rect 376018 22788 376024 22840
rect 376076 22828 376082 22840
rect 452746 22828 452752 22840
rect 376076 22800 452752 22828
rect 376076 22788 376082 22800
rect 452746 22788 452752 22800
rect 452804 22788 452810 22840
rect 238018 22720 238024 22772
rect 238076 22760 238082 22772
rect 394694 22760 394700 22772
rect 238076 22732 394700 22760
rect 238076 22720 238082 22732
rect 394694 22720 394700 22732
rect 394752 22720 394758 22772
rect 224770 21428 224776 21480
rect 224828 21468 224834 21480
rect 345014 21468 345020 21480
rect 224828 21440 345020 21468
rect 224828 21428 224834 21440
rect 345014 21428 345020 21440
rect 345072 21428 345078 21480
rect 238018 21360 238024 21412
rect 238076 21400 238082 21412
rect 423674 21400 423680 21412
rect 238076 21372 423680 21400
rect 238076 21360 238082 21372
rect 423674 21360 423680 21372
rect 423732 21360 423738 21412
rect 519630 20612 519636 20664
rect 519688 20652 519694 20664
rect 579982 20652 579988 20664
rect 519688 20624 579988 20652
rect 519688 20612 519694 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 228358 20000 228364 20052
rect 228416 20040 228422 20052
rect 334066 20040 334072 20052
rect 228416 20012 334072 20040
rect 228416 20000 228422 20012
rect 334066 20000 334072 20012
rect 334124 20000 334130 20052
rect 374638 20000 374644 20052
rect 374696 20040 374702 20052
rect 454034 20040 454040 20052
rect 374696 20012 454040 20040
rect 374696 20000 374702 20012
rect 454034 20000 454040 20012
rect 454092 20000 454098 20052
rect 59262 19932 59268 19984
rect 59320 19972 59326 19984
rect 85574 19972 85580 19984
rect 59320 19944 85580 19972
rect 59320 19932 59326 19944
rect 85574 19932 85580 19944
rect 85632 19932 85638 19984
rect 224770 19932 224776 19984
rect 224828 19972 224834 19984
rect 410518 19972 410524 19984
rect 224828 19944 410524 19972
rect 224828 19932 224834 19944
rect 410518 19932 410524 19944
rect 410576 19932 410582 19984
rect 220078 18640 220084 18692
rect 220136 18680 220142 18692
rect 324406 18680 324412 18692
rect 220136 18652 324412 18680
rect 220136 18640 220142 18652
rect 324406 18640 324412 18652
rect 324464 18640 324470 18692
rect 68370 18572 68376 18624
rect 68428 18612 68434 18624
rect 143534 18612 143540 18624
rect 68428 18584 143540 18612
rect 68428 18572 68434 18584
rect 143534 18572 143540 18584
rect 143592 18572 143598 18624
rect 220630 18572 220636 18624
rect 220688 18612 220694 18624
rect 421558 18612 421564 18624
rect 220688 18584 421564 18612
rect 220688 18572 220694 18584
rect 421558 18572 421564 18584
rect 421616 18572 421622 18624
rect 358078 17484 358084 17536
rect 358136 17524 358142 17536
rect 409966 17524 409972 17536
rect 358136 17496 409972 17524
rect 358136 17484 358142 17496
rect 409966 17484 409972 17496
rect 410024 17484 410030 17536
rect 216490 17416 216496 17468
rect 216548 17456 216554 17468
rect 313366 17456 313372 17468
rect 216548 17428 313372 17456
rect 216548 17416 216554 17428
rect 313366 17416 313372 17428
rect 313424 17416 313430 17468
rect 358170 17416 358176 17468
rect 358228 17456 358234 17468
rect 448606 17456 448612 17468
rect 358228 17428 448612 17456
rect 358228 17416 358234 17428
rect 448606 17416 448612 17428
rect 448664 17416 448670 17468
rect 294598 17348 294604 17400
rect 294656 17388 294662 17400
rect 438854 17388 438860 17400
rect 294656 17360 438860 17388
rect 294656 17348 294662 17360
rect 438854 17348 438860 17360
rect 438912 17348 438918 17400
rect 269758 17280 269764 17332
rect 269816 17320 269822 17332
rect 430574 17320 430580 17332
rect 269816 17292 430580 17320
rect 269816 17280 269822 17292
rect 430574 17280 430580 17292
rect 430632 17280 430638 17332
rect 32398 17212 32404 17264
rect 32456 17252 32462 17264
rect 78674 17252 78680 17264
rect 32456 17224 78680 17252
rect 32456 17212 32462 17224
rect 78674 17212 78680 17224
rect 78732 17212 78738 17264
rect 143442 17212 143448 17264
rect 143500 17252 143506 17264
rect 392578 17252 392584 17264
rect 143500 17224 392584 17252
rect 143500 17212 143506 17224
rect 392578 17212 392584 17224
rect 392636 17212 392642 17264
rect 211062 16260 211068 16312
rect 211120 16300 211126 16312
rect 295610 16300 295616 16312
rect 211120 16272 295616 16300
rect 211120 16260 211126 16272
rect 295610 16260 295616 16272
rect 295668 16260 295674 16312
rect 377950 16192 377956 16244
rect 378008 16232 378014 16244
rect 468478 16232 468484 16244
rect 378008 16204 468484 16232
rect 378008 16192 378014 16204
rect 468478 16192 468484 16204
rect 468536 16192 468542 16244
rect 180058 16124 180064 16176
rect 180116 16164 180122 16176
rect 295426 16164 295432 16176
rect 180116 16136 295432 16164
rect 180116 16124 180122 16136
rect 295426 16124 295432 16136
rect 295484 16124 295490 16176
rect 323578 16124 323584 16176
rect 323636 16164 323642 16176
rect 447134 16164 447140 16176
rect 323636 16136 447140 16164
rect 323636 16124 323642 16136
rect 447134 16124 447140 16136
rect 447192 16124 447198 16176
rect 291838 16056 291844 16108
rect 291896 16096 291902 16108
rect 436094 16096 436100 16108
rect 291896 16068 436100 16096
rect 291896 16056 291902 16068
rect 436094 16056 436100 16068
rect 436152 16056 436158 16108
rect 240870 15988 240876 16040
rect 240928 16028 240934 16040
rect 425054 16028 425060 16040
rect 240928 16000 425060 16028
rect 240928 15988 240934 16000
rect 425054 15988 425060 16000
rect 425112 15988 425118 16040
rect 220078 15920 220084 15972
rect 220136 15960 220142 15972
rect 420914 15960 420920 15972
rect 220136 15932 420920 15960
rect 220136 15920 220142 15932
rect 420914 15920 420920 15932
rect 420972 15920 420978 15972
rect 52362 15852 52368 15904
rect 52420 15892 52426 15904
rect 68278 15892 68284 15904
rect 52420 15864 68284 15892
rect 52420 15852 52426 15864
rect 68278 15852 68284 15864
rect 68336 15852 68342 15904
rect 139302 15852 139308 15904
rect 139360 15892 139366 15904
rect 400858 15892 400864 15904
rect 139360 15864 400864 15892
rect 139360 15852 139366 15864
rect 400858 15852 400864 15864
rect 400916 15852 400922 15904
rect 259270 14900 259276 14952
rect 259328 14940 259334 14952
rect 316034 14940 316040 14952
rect 259328 14912 316040 14940
rect 259328 14900 259334 14912
rect 316034 14900 316040 14912
rect 316092 14900 316098 14952
rect 169570 14832 169576 14884
rect 169628 14872 169634 14884
rect 289078 14872 289084 14884
rect 169628 14844 289084 14872
rect 169628 14832 169634 14844
rect 289078 14832 289084 14844
rect 289136 14832 289142 14884
rect 377398 14832 377404 14884
rect 377456 14872 377462 14884
rect 452654 14872 452660 14884
rect 377456 14844 452660 14872
rect 377456 14832 377462 14844
rect 452654 14832 452660 14844
rect 452712 14832 452718 14884
rect 144730 14764 144736 14816
rect 144788 14804 144794 14816
rect 287054 14804 287060 14816
rect 144788 14776 287060 14804
rect 144788 14764 144794 14776
rect 287054 14764 287060 14776
rect 287112 14764 287118 14816
rect 287790 14764 287796 14816
rect 287848 14804 287854 14816
rect 434714 14804 434720 14816
rect 287848 14776 434720 14804
rect 287848 14764 287854 14776
rect 434714 14764 434720 14776
rect 434772 14764 434778 14816
rect 137646 14696 137652 14748
rect 137704 14736 137710 14748
rect 285674 14736 285680 14748
rect 137704 14708 285680 14736
rect 137704 14696 137710 14708
rect 285674 14696 285680 14708
rect 285732 14696 285738 14748
rect 292482 14696 292488 14748
rect 292540 14736 292546 14748
rect 439498 14736 439504 14748
rect 292540 14708 439504 14736
rect 292540 14696 292546 14708
rect 439498 14696 439504 14708
rect 439556 14696 439562 14748
rect 240778 14628 240784 14680
rect 240836 14668 240842 14680
rect 398834 14668 398840 14680
rect 240836 14640 398840 14668
rect 240836 14628 240842 14640
rect 398834 14628 398840 14640
rect 398892 14628 398898 14680
rect 246298 14560 246304 14612
rect 246356 14600 246362 14612
rect 406010 14600 406016 14612
rect 246356 14572 406016 14600
rect 246356 14560 246362 14572
rect 406010 14560 406016 14572
rect 406068 14560 406074 14612
rect 246390 14492 246396 14544
rect 246448 14532 246454 14544
rect 427814 14532 427820 14544
rect 246448 14504 427820 14532
rect 246448 14492 246454 14504
rect 427814 14492 427820 14504
rect 427872 14492 427878 14544
rect 54938 14424 54944 14476
rect 54996 14464 55002 14476
rect 65610 14464 65616 14476
rect 54996 14436 65616 14464
rect 54996 14424 55002 14436
rect 65610 14424 65616 14436
rect 65668 14424 65674 14476
rect 259362 14424 259368 14476
rect 259420 14464 259426 14476
rect 483658 14464 483664 14476
rect 259420 14436 483664 14464
rect 259420 14424 259426 14436
rect 483658 14424 483664 14436
rect 483716 14424 483722 14476
rect 268838 13676 268844 13728
rect 268896 13716 268902 13728
rect 316678 13716 316684 13728
rect 268896 13688 316684 13716
rect 268896 13676 268902 13688
rect 316678 13676 316684 13688
rect 316736 13676 316742 13728
rect 216582 13608 216588 13660
rect 216640 13648 216646 13660
rect 316034 13648 316040 13660
rect 216640 13620 316040 13648
rect 216640 13608 216646 13620
rect 316034 13608 316040 13620
rect 316092 13608 316098 13660
rect 220722 13540 220728 13592
rect 220780 13580 220786 13592
rect 331582 13580 331588 13592
rect 220780 13552 331588 13580
rect 220780 13540 220786 13552
rect 331582 13540 331588 13552
rect 331640 13540 331646 13592
rect 379422 13540 379428 13592
rect 379480 13580 379486 13592
rect 471238 13580 471244 13592
rect 379480 13552 471244 13580
rect 379480 13540 379486 13552
rect 471238 13540 471244 13552
rect 471296 13540 471302 13592
rect 224862 13472 224868 13524
rect 224920 13512 224926 13524
rect 349246 13512 349252 13524
rect 224920 13484 349252 13512
rect 224920 13472 224926 13484
rect 349246 13472 349252 13484
rect 349304 13472 349310 13524
rect 353938 13472 353944 13524
rect 353996 13512 354002 13524
rect 448514 13512 448520 13524
rect 353996 13484 448520 13512
rect 353996 13472 354002 13484
rect 448514 13472 448520 13484
rect 448572 13472 448578 13524
rect 180702 13404 180708 13456
rect 180760 13444 180766 13456
rect 295978 13444 295984 13456
rect 180760 13416 295984 13444
rect 180760 13404 180766 13416
rect 295978 13404 295984 13416
rect 296036 13404 296042 13456
rect 316770 13404 316776 13456
rect 316828 13444 316834 13456
rect 442994 13444 443000 13456
rect 316828 13416 443000 13444
rect 316828 13404 316834 13416
rect 442994 13404 443000 13416
rect 443052 13404 443058 13456
rect 227530 13336 227536 13388
rect 227588 13376 227594 13388
rect 356330 13376 356336 13388
rect 227588 13348 356336 13376
rect 227588 13336 227594 13348
rect 356330 13336 356336 13348
rect 356388 13336 356394 13388
rect 378042 13336 378048 13388
rect 378100 13376 378106 13388
rect 497458 13376 497464 13388
rect 378100 13348 497464 13376
rect 378100 13336 378106 13348
rect 497458 13336 497464 13348
rect 497516 13336 497522 13388
rect 281258 13268 281264 13320
rect 281316 13308 281322 13320
rect 431218 13308 431224 13320
rect 281316 13280 431224 13308
rect 281316 13268 281322 13280
rect 431218 13268 431224 13280
rect 431276 13268 431282 13320
rect 234522 13200 234528 13252
rect 234580 13240 234586 13252
rect 387794 13240 387800 13252
rect 234580 13212 387800 13240
rect 234580 13200 234586 13212
rect 387794 13200 387800 13212
rect 387852 13200 387858 13252
rect 264330 13132 264336 13184
rect 264388 13172 264394 13184
rect 431954 13172 431960 13184
rect 264388 13144 431960 13172
rect 264388 13132 264394 13144
rect 431954 13132 431960 13144
rect 432012 13132 432018 13184
rect 17862 13064 17868 13116
rect 17920 13104 17926 13116
rect 75914 13104 75920 13116
rect 17920 13076 75920 13104
rect 17920 13064 17926 13076
rect 75914 13064 75920 13076
rect 75972 13064 75978 13116
rect 76558 13064 76564 13116
rect 76616 13104 76622 13116
rect 147766 13104 147772 13116
rect 76616 13076 147772 13104
rect 76616 13064 76622 13076
rect 147766 13064 147772 13076
rect 147824 13064 147830 13116
rect 202138 13064 202144 13116
rect 202196 13104 202202 13116
rect 214466 13104 214472 13116
rect 202196 13076 214472 13104
rect 202196 13064 202202 13076
rect 214466 13064 214472 13076
rect 214524 13064 214530 13116
rect 264882 13064 264888 13116
rect 264940 13104 264946 13116
rect 504358 13104 504364 13116
rect 264940 13076 504364 13104
rect 264940 13064 264946 13076
rect 504358 13064 504364 13076
rect 504416 13064 504422 13116
rect 209682 12384 209688 12436
rect 209740 12424 209746 12436
rect 288986 12424 288992 12436
rect 209740 12396 288992 12424
rect 209740 12384 209746 12396
rect 288986 12384 288992 12396
rect 289044 12384 289050 12436
rect 213822 12316 213828 12368
rect 213880 12356 213886 12368
rect 303154 12356 303160 12368
rect 213880 12328 303160 12356
rect 213880 12316 213886 12328
rect 303154 12316 303160 12328
rect 303212 12316 303218 12368
rect 378778 12316 378784 12368
rect 378836 12356 378842 12368
rect 403618 12356 403624 12368
rect 378836 12328 403624 12356
rect 378836 12316 378842 12328
rect 403618 12316 403624 12328
rect 403676 12316 403682 12368
rect 215202 12248 215208 12300
rect 215260 12288 215266 12300
rect 309778 12288 309784 12300
rect 215260 12260 309784 12288
rect 215260 12248 215266 12260
rect 309778 12248 309784 12260
rect 309836 12248 309842 12300
rect 354582 12248 354588 12300
rect 354640 12288 354646 12300
rect 407114 12288 407120 12300
rect 354640 12260 407120 12288
rect 354640 12248 354646 12260
rect 407114 12248 407120 12260
rect 407172 12248 407178 12300
rect 223482 12180 223488 12232
rect 223540 12220 223546 12232
rect 340874 12220 340880 12232
rect 223540 12192 340880 12220
rect 223540 12180 223546 12192
rect 340874 12180 340880 12192
rect 340932 12180 340938 12232
rect 375282 12180 375288 12232
rect 375340 12220 375346 12232
rect 484762 12220 484768 12232
rect 375340 12192 484768 12220
rect 375340 12180 375346 12192
rect 484762 12180 484768 12192
rect 484820 12180 484826 12232
rect 217962 12112 217968 12164
rect 218020 12152 218026 12164
rect 320450 12152 320456 12164
rect 218020 12124 320456 12152
rect 218020 12112 218026 12124
rect 320450 12112 320456 12124
rect 320508 12112 320514 12164
rect 322290 12112 322296 12164
rect 322348 12152 322354 12164
rect 445846 12152 445852 12164
rect 322348 12124 445852 12152
rect 322348 12112 322354 12124
rect 445846 12112 445852 12124
rect 445904 12112 445910 12164
rect 227622 12044 227628 12096
rect 227680 12084 227686 12096
rect 359458 12084 359464 12096
rect 227680 12056 359464 12084
rect 227680 12044 227686 12056
rect 359458 12044 359464 12056
rect 359516 12044 359522 12096
rect 376662 12044 376668 12096
rect 376720 12084 376726 12096
rect 490558 12084 490564 12096
rect 376720 12056 490564 12084
rect 376720 12044 376726 12056
rect 490558 12044 490564 12056
rect 490616 12044 490622 12096
rect 285582 11976 285588 12028
rect 285640 12016 285646 12028
rect 436738 12016 436744 12028
rect 285640 11988 436744 12016
rect 285640 11976 285646 11988
rect 436738 11976 436744 11988
rect 436796 11976 436802 12028
rect 238662 11908 238668 11960
rect 238720 11948 238726 11960
rect 402514 11948 402520 11960
rect 238720 11920 402520 11948
rect 238720 11908 238726 11920
rect 402514 11908 402520 11920
rect 402572 11908 402578 11960
rect 260650 11840 260656 11892
rect 260708 11880 260714 11892
rect 489270 11880 489276 11892
rect 260708 11852 489276 11880
rect 260708 11840 260714 11852
rect 489270 11840 489276 11852
rect 489328 11840 489334 11892
rect 57330 11772 57336 11824
rect 57388 11812 57394 11824
rect 142154 11812 142160 11824
rect 57388 11784 142160 11812
rect 57388 11772 57394 11784
rect 142154 11772 142160 11784
rect 142212 11772 142218 11824
rect 263410 11772 263416 11824
rect 263468 11812 263474 11824
rect 501322 11812 501328 11824
rect 263468 11784 501328 11812
rect 263468 11772 263474 11784
rect 501322 11772 501328 11784
rect 501380 11772 501386 11824
rect 136450 11704 136456 11756
rect 136508 11744 136514 11756
rect 381538 11744 381544 11756
rect 136508 11716 381544 11744
rect 136508 11704 136514 11716
rect 381538 11704 381544 11716
rect 381596 11704 381602 11756
rect 192938 10956 192944 11008
rect 192996 10996 193002 11008
rect 414014 10996 414020 11008
rect 192996 10968 414020 10996
rect 192996 10956 193002 10968
rect 414014 10956 414020 10968
rect 414072 10956 414078 11008
rect 188982 10888 188988 10940
rect 189040 10928 189046 10940
rect 414106 10928 414112 10940
rect 189040 10900 414112 10928
rect 189040 10888 189046 10900
rect 414106 10888 414112 10900
rect 414164 10888 414170 10940
rect 186222 10820 186228 10872
rect 186280 10860 186286 10872
rect 412634 10860 412640 10872
rect 186280 10832 412640 10860
rect 186280 10820 186286 10832
rect 412634 10820 412640 10832
rect 412692 10820 412698 10872
rect 182082 10752 182088 10804
rect 182140 10792 182146 10804
rect 411254 10792 411260 10804
rect 182140 10764 411260 10792
rect 182140 10752 182146 10764
rect 411254 10752 411260 10764
rect 411312 10752 411318 10804
rect 177850 10684 177856 10736
rect 177908 10724 177914 10736
rect 411346 10724 411352 10736
rect 177908 10696 411352 10724
rect 177908 10684 177914 10696
rect 411346 10684 411352 10696
rect 411404 10684 411410 10736
rect 175182 10616 175188 10668
rect 175240 10656 175246 10668
rect 409874 10656 409880 10668
rect 175240 10628 409880 10656
rect 175240 10616 175246 10628
rect 409874 10616 409880 10628
rect 409932 10616 409938 10668
rect 170766 10548 170772 10600
rect 170824 10588 170830 10600
rect 408586 10588 408592 10600
rect 170824 10560 408592 10588
rect 170824 10548 170830 10560
rect 408586 10548 408592 10560
rect 408644 10548 408650 10600
rect 168282 10480 168288 10532
rect 168340 10520 168346 10532
rect 408494 10520 408500 10532
rect 168340 10492 408500 10520
rect 168340 10480 168346 10492
rect 408494 10480 408500 10492
rect 408552 10480 408558 10532
rect 164142 10412 164148 10464
rect 164200 10452 164206 10464
rect 407206 10452 407212 10464
rect 164200 10424 407212 10452
rect 164200 10412 164206 10424
rect 407206 10412 407212 10424
rect 407264 10412 407270 10464
rect 131758 10344 131764 10396
rect 131816 10384 131822 10396
rect 399018 10384 399024 10396
rect 131816 10356 399024 10384
rect 131816 10344 131822 10356
rect 399018 10344 399024 10356
rect 399076 10344 399082 10396
rect 66162 10276 66168 10328
rect 66220 10316 66226 10328
rect 86954 10316 86960 10328
rect 66220 10288 86960 10316
rect 66220 10276 66226 10288
rect 86954 10276 86960 10288
rect 87012 10276 87018 10328
rect 128170 10276 128176 10328
rect 128228 10316 128234 10328
rect 398926 10316 398932 10328
rect 128228 10288 398932 10316
rect 128228 10276 128234 10288
rect 398926 10276 398932 10288
rect 398984 10276 398990 10328
rect 418798 10276 418804 10328
rect 418856 10316 418862 10328
rect 506474 10316 506480 10328
rect 418856 10288 506480 10316
rect 418856 10276 418862 10288
rect 506474 10276 506480 10288
rect 506532 10276 506538 10328
rect 195606 10208 195612 10260
rect 195664 10248 195670 10260
rect 415394 10248 415400 10260
rect 195664 10220 415400 10248
rect 195664 10208 195670 10220
rect 415394 10208 415400 10220
rect 415452 10208 415458 10260
rect 199930 10140 199936 10192
rect 199988 10180 199994 10192
rect 416866 10180 416872 10192
rect 199988 10152 416872 10180
rect 199988 10140 199994 10152
rect 416866 10140 416872 10152
rect 416924 10140 416930 10192
rect 202690 10072 202696 10124
rect 202748 10112 202754 10124
rect 416774 10112 416780 10124
rect 202748 10084 416780 10112
rect 202748 10072 202754 10084
rect 416774 10072 416780 10084
rect 416832 10072 416838 10124
rect 206738 10004 206744 10056
rect 206796 10044 206802 10056
rect 418154 10044 418160 10056
rect 206796 10016 418160 10044
rect 206796 10004 206802 10016
rect 418154 10004 418160 10016
rect 418212 10004 418218 10056
rect 211062 9936 211068 9988
rect 211120 9976 211126 9988
rect 419626 9976 419632 9988
rect 211120 9948 419632 9976
rect 211120 9936 211126 9948
rect 419626 9936 419632 9948
rect 419684 9936 419690 9988
rect 213822 9868 213828 9920
rect 213880 9908 213886 9920
rect 419534 9908 419540 9920
rect 213880 9880 419540 9908
rect 213880 9868 213886 9880
rect 419534 9868 419540 9880
rect 419592 9868 419598 9920
rect 277118 9800 277124 9852
rect 277176 9840 277182 9852
rect 320266 9840 320272 9852
rect 277176 9812 320272 9840
rect 277176 9800 277182 9812
rect 320266 9800 320272 9812
rect 320324 9800 320330 9852
rect 279510 9732 279516 9784
rect 279568 9772 279574 9784
rect 321554 9772 321560 9784
rect 279568 9744 321560 9772
rect 279568 9732 279574 9744
rect 321554 9732 321560 9744
rect 321612 9732 321618 9784
rect 222746 9596 222752 9648
rect 222804 9636 222810 9648
rect 306466 9636 306472 9648
rect 222804 9608 306472 9636
rect 222804 9596 222810 9608
rect 306466 9596 306472 9608
rect 306524 9596 306530 9648
rect 364242 9596 364248 9648
rect 364300 9636 364306 9648
rect 442626 9636 442632 9648
rect 364300 9608 442632 9636
rect 364300 9596 364306 9608
rect 442626 9596 442632 9608
rect 442684 9596 442690 9648
rect 219250 9528 219256 9580
rect 219308 9568 219314 9580
rect 306374 9568 306380 9580
rect 219308 9540 306380 9568
rect 219308 9528 219314 9540
rect 306374 9528 306380 9540
rect 306432 9528 306438 9580
rect 365530 9528 365536 9580
rect 365588 9568 365594 9580
rect 446214 9568 446220 9580
rect 365588 9540 446220 9568
rect 365588 9528 365594 9540
rect 446214 9528 446220 9540
rect 446272 9528 446278 9580
rect 215662 9460 215668 9512
rect 215720 9500 215726 9512
rect 304994 9500 305000 9512
rect 215720 9472 305000 9500
rect 215720 9460 215726 9472
rect 304994 9460 305000 9472
rect 305052 9460 305058 9512
rect 365622 9460 365628 9512
rect 365680 9500 365686 9512
rect 449802 9500 449808 9512
rect 365680 9472 449808 9500
rect 365680 9460 365686 9472
rect 449802 9460 449808 9472
rect 449860 9460 449866 9512
rect 212166 9392 212172 9444
rect 212224 9432 212230 9444
rect 303614 9432 303620 9444
rect 212224 9404 303620 9432
rect 212224 9392 212230 9404
rect 303614 9392 303620 9404
rect 303672 9392 303678 9444
rect 367002 9392 367008 9444
rect 367060 9432 367066 9444
rect 453298 9432 453304 9444
rect 367060 9404 453304 9432
rect 367060 9392 367066 9404
rect 453298 9392 453304 9404
rect 453356 9392 453362 9444
rect 208578 9324 208584 9376
rect 208636 9364 208642 9376
rect 303706 9364 303712 9376
rect 208636 9336 303712 9364
rect 208636 9324 208642 9336
rect 303706 9324 303712 9336
rect 303764 9324 303770 9376
rect 368382 9324 368388 9376
rect 368440 9364 368446 9376
rect 456886 9364 456892 9376
rect 368440 9336 456892 9364
rect 368440 9324 368446 9336
rect 456886 9324 456892 9336
rect 456944 9324 456950 9376
rect 205082 9256 205088 9308
rect 205140 9296 205146 9308
rect 302418 9296 302424 9308
rect 205140 9268 302424 9296
rect 205140 9256 205146 9268
rect 302418 9256 302424 9268
rect 302476 9256 302482 9308
rect 368290 9256 368296 9308
rect 368348 9296 368354 9308
rect 460382 9296 460388 9308
rect 368348 9268 460388 9296
rect 368348 9256 368354 9268
rect 460382 9256 460388 9268
rect 460440 9256 460446 9308
rect 201494 9188 201500 9240
rect 201552 9228 201558 9240
rect 302326 9228 302332 9240
rect 201552 9200 302332 9228
rect 201552 9188 201558 9200
rect 302326 9188 302332 9200
rect 302384 9188 302390 9240
rect 369762 9188 369768 9240
rect 369820 9228 369826 9240
rect 463970 9228 463976 9240
rect 369820 9200 463976 9228
rect 369820 9188 369826 9200
rect 463970 9188 463976 9200
rect 464028 9188 464034 9240
rect 197906 9120 197912 9172
rect 197964 9160 197970 9172
rect 300854 9160 300860 9172
rect 197964 9132 300860 9160
rect 197964 9120 197970 9132
rect 300854 9120 300860 9132
rect 300912 9120 300918 9172
rect 371142 9120 371148 9172
rect 371200 9160 371206 9172
rect 467466 9160 467472 9172
rect 371200 9132 467472 9160
rect 371200 9120 371206 9132
rect 467466 9120 467472 9132
rect 467524 9120 467530 9172
rect 194410 9052 194416 9104
rect 194468 9092 194474 9104
rect 299474 9092 299480 9104
rect 194468 9064 299480 9092
rect 194468 9052 194474 9064
rect 299474 9052 299480 9064
rect 299532 9052 299538 9104
rect 325602 9052 325608 9104
rect 325660 9092 325666 9104
rect 331858 9092 331864 9104
rect 325660 9064 331864 9092
rect 325660 9052 325666 9064
rect 331858 9052 331864 9064
rect 331916 9052 331922 9104
rect 371050 9052 371056 9104
rect 371108 9092 371114 9104
rect 471054 9092 471060 9104
rect 371108 9064 471060 9092
rect 371108 9052 371114 9064
rect 471054 9052 471060 9064
rect 471112 9052 471118 9104
rect 69658 9024 69664 9036
rect 64846 8996 69664 9024
rect 47854 8916 47860 8968
rect 47912 8956 47918 8968
rect 64846 8956 64874 8996
rect 69658 8984 69664 8996
rect 69716 8984 69722 9036
rect 134150 8984 134156 9036
rect 134208 9024 134214 9036
rect 284294 9024 284300 9036
rect 134208 8996 284300 9024
rect 134208 8984 134214 8996
rect 284294 8984 284300 8996
rect 284352 8984 284358 9036
rect 322198 8984 322204 9036
rect 322256 9024 322262 9036
rect 338666 9024 338672 9036
rect 322256 8996 338672 9024
rect 322256 8984 322262 8996
rect 338666 8984 338672 8996
rect 338724 8984 338730 9036
rect 340138 8984 340144 9036
rect 340196 9024 340202 9036
rect 352834 9024 352840 9036
rect 340196 8996 352840 9024
rect 340196 8984 340202 8996
rect 352834 8984 352840 8996
rect 352892 8984 352898 9036
rect 372522 8984 372528 9036
rect 372580 9024 372586 9036
rect 474550 9024 474556 9036
rect 372580 8996 474556 9024
rect 372580 8984 372586 8996
rect 474550 8984 474556 8996
rect 474608 8984 474614 9036
rect 47912 8928 64874 8956
rect 47912 8916 47918 8928
rect 69106 8916 69112 8968
rect 69164 8956 69170 8968
rect 88334 8956 88340 8968
rect 69164 8928 88340 8956
rect 69164 8916 69170 8928
rect 88334 8916 88340 8928
rect 88392 8916 88398 8968
rect 105722 8916 105728 8968
rect 105780 8956 105786 8968
rect 124858 8956 124864 8968
rect 105780 8928 124864 8956
rect 105780 8916 105786 8928
rect 124858 8916 124864 8928
rect 124916 8916 124922 8968
rect 130562 8916 130568 8968
rect 130620 8956 130626 8968
rect 283006 8956 283012 8968
rect 130620 8928 283012 8956
rect 130620 8916 130626 8928
rect 283006 8916 283012 8928
rect 283064 8916 283070 8968
rect 312630 8916 312636 8968
rect 312688 8956 312694 8968
rect 353846 8956 353852 8968
rect 312688 8928 353852 8956
rect 312688 8916 312694 8928
rect 353846 8916 353852 8928
rect 353904 8916 353910 8968
rect 373902 8916 373908 8968
rect 373960 8956 373966 8968
rect 478138 8956 478144 8968
rect 373960 8928 478144 8956
rect 373960 8916 373966 8928
rect 478138 8916 478144 8928
rect 478196 8916 478202 8968
rect 226334 8848 226340 8900
rect 226392 8888 226398 8900
rect 307754 8888 307760 8900
rect 226392 8860 307760 8888
rect 226392 8848 226398 8860
rect 307754 8848 307760 8860
rect 307812 8848 307818 8900
rect 362770 8848 362776 8900
rect 362828 8888 362834 8900
rect 439130 8888 439136 8900
rect 362828 8860 439136 8888
rect 362828 8848 362834 8860
rect 439130 8848 439136 8860
rect 439188 8848 439194 8900
rect 229830 8780 229836 8832
rect 229888 8820 229894 8832
rect 309226 8820 309232 8832
rect 229888 8792 309232 8820
rect 229888 8780 229894 8792
rect 309226 8780 309232 8792
rect 309284 8780 309290 8832
rect 362862 8780 362868 8832
rect 362920 8820 362926 8832
rect 435542 8820 435548 8832
rect 362920 8792 435548 8820
rect 362920 8780 362926 8792
rect 435542 8780 435548 8792
rect 435600 8780 435606 8832
rect 233418 8712 233424 8764
rect 233476 8752 233482 8764
rect 309318 8752 309324 8764
rect 233476 8724 309324 8752
rect 233476 8712 233482 8724
rect 309318 8712 309324 8724
rect 309376 8712 309382 8764
rect 361482 8712 361488 8764
rect 361540 8752 361546 8764
rect 432046 8752 432052 8764
rect 361540 8724 432052 8752
rect 361540 8712 361546 8724
rect 432046 8712 432052 8724
rect 432104 8712 432110 8764
rect 237006 8644 237012 8696
rect 237064 8684 237070 8696
rect 310514 8684 310520 8696
rect 237064 8656 310520 8684
rect 237064 8644 237070 8656
rect 310514 8644 310520 8656
rect 310572 8644 310578 8696
rect 360010 8644 360016 8696
rect 360068 8684 360074 8696
rect 428458 8684 428464 8696
rect 360068 8656 428464 8684
rect 360068 8644 360074 8656
rect 428458 8644 428464 8656
rect 428516 8644 428522 8696
rect 240502 8576 240508 8628
rect 240560 8616 240566 8628
rect 311894 8616 311900 8628
rect 240560 8588 311900 8616
rect 240560 8576 240566 8588
rect 311894 8576 311900 8588
rect 311952 8576 311958 8628
rect 360102 8576 360108 8628
rect 360160 8616 360166 8628
rect 424962 8616 424968 8628
rect 360160 8588 424968 8616
rect 360160 8576 360166 8588
rect 424962 8576 424968 8588
rect 425020 8576 425026 8628
rect 244090 8508 244096 8560
rect 244148 8548 244154 8560
rect 311986 8548 311992 8560
rect 244148 8520 311992 8548
rect 244148 8508 244154 8520
rect 311986 8508 311992 8520
rect 312044 8508 312050 8560
rect 358722 8508 358728 8560
rect 358780 8548 358786 8560
rect 421374 8548 421380 8560
rect 358780 8520 421380 8548
rect 358780 8508 358786 8520
rect 421374 8508 421380 8520
rect 421432 8508 421438 8560
rect 247586 8440 247592 8492
rect 247644 8480 247650 8492
rect 313274 8480 313280 8492
rect 247644 8452 313280 8480
rect 247644 8440 247650 8452
rect 313274 8440 313280 8452
rect 313332 8440 313338 8492
rect 357342 8440 357348 8492
rect 357400 8480 357406 8492
rect 417878 8480 417884 8492
rect 357400 8452 417884 8480
rect 357400 8440 357406 8452
rect 417878 8440 417884 8452
rect 417936 8440 417942 8492
rect 251174 8372 251180 8424
rect 251232 8412 251238 8424
rect 314746 8412 314752 8424
rect 251232 8384 314752 8412
rect 251232 8372 251238 8384
rect 314746 8372 314752 8384
rect 314804 8372 314810 8424
rect 357250 8372 357256 8424
rect 357308 8412 357314 8424
rect 414290 8412 414296 8424
rect 357308 8384 414296 8412
rect 357308 8372 357314 8384
rect 414290 8372 414296 8384
rect 414348 8372 414354 8424
rect 305638 8304 305644 8356
rect 305696 8344 305702 8356
rect 306742 8344 306748 8356
rect 305696 8316 306748 8344
rect 305696 8304 305702 8316
rect 306742 8304 306748 8316
rect 306800 8304 306806 8356
rect 52546 8236 52552 8288
rect 52604 8276 52610 8288
rect 54478 8276 54484 8288
rect 52604 8248 54484 8276
rect 52604 8236 52610 8248
rect 54478 8236 54484 8248
rect 54536 8236 54542 8288
rect 248230 8236 248236 8288
rect 248288 8276 248294 8288
rect 441246 8276 441252 8288
rect 248288 8248 441252 8276
rect 248288 8236 248294 8248
rect 441246 8236 441252 8248
rect 441304 8236 441310 8288
rect 249702 8168 249708 8220
rect 249760 8208 249766 8220
rect 445018 8208 445024 8220
rect 249760 8180 445024 8208
rect 249760 8168 249766 8180
rect 445018 8168 445024 8180
rect 445076 8168 445082 8220
rect 250990 8100 250996 8152
rect 251048 8140 251054 8152
rect 448606 8140 448612 8152
rect 251048 8112 448612 8140
rect 251048 8100 251054 8112
rect 448606 8100 448612 8112
rect 448664 8100 448670 8152
rect 450538 8100 450544 8152
rect 450596 8140 450602 8152
rect 480530 8140 480536 8152
rect 450596 8112 480536 8140
rect 450596 8100 450602 8112
rect 480530 8100 480536 8112
rect 480588 8100 480594 8152
rect 251082 8032 251088 8084
rect 251140 8072 251146 8084
rect 452102 8072 452108 8084
rect 251140 8044 452108 8072
rect 251140 8032 251146 8044
rect 452102 8032 452108 8044
rect 452160 8032 452166 8084
rect 252462 7964 252468 8016
rect 252520 8004 252526 8016
rect 455690 8004 455696 8016
rect 252520 7976 455696 8004
rect 252520 7964 252526 7976
rect 455690 7964 455696 7976
rect 455748 7964 455754 8016
rect 253750 7896 253756 7948
rect 253808 7936 253814 7948
rect 459186 7936 459192 7948
rect 253808 7908 459192 7936
rect 253808 7896 253814 7908
rect 459186 7896 459192 7908
rect 459244 7896 459250 7948
rect 253842 7828 253848 7880
rect 253900 7868 253906 7880
rect 462774 7868 462780 7880
rect 253900 7840 462780 7868
rect 253900 7828 253906 7840
rect 462774 7828 462780 7840
rect 462832 7828 462838 7880
rect 255222 7760 255228 7812
rect 255280 7800 255286 7812
rect 466270 7800 466276 7812
rect 255280 7772 466276 7800
rect 255280 7760 255286 7772
rect 466270 7760 466276 7772
rect 466328 7760 466334 7812
rect 256602 7692 256608 7744
rect 256660 7732 256666 7744
rect 469858 7732 469864 7744
rect 256660 7704 469864 7732
rect 256660 7692 256666 7704
rect 469858 7692 469864 7704
rect 469916 7692 469922 7744
rect 70302 7624 70308 7676
rect 70360 7664 70366 7676
rect 118694 7664 118700 7676
rect 70360 7636 118700 7664
rect 70360 7624 70366 7636
rect 118694 7624 118700 7636
rect 118752 7624 118758 7676
rect 256510 7624 256516 7676
rect 256568 7664 256574 7676
rect 473446 7664 473452 7676
rect 256568 7636 473452 7664
rect 256568 7624 256574 7636
rect 473446 7624 473452 7636
rect 473504 7624 473510 7676
rect 42978 7556 42984 7608
rect 43036 7596 43042 7608
rect 110414 7596 110420 7608
rect 43036 7568 110420 7596
rect 43036 7556 43042 7568
rect 110414 7556 110420 7568
rect 110472 7556 110478 7608
rect 119890 7556 119896 7608
rect 119948 7596 119954 7608
rect 128998 7596 129004 7608
rect 119948 7568 129004 7596
rect 119948 7556 119954 7568
rect 128998 7556 129004 7568
rect 129056 7556 129062 7608
rect 257982 7556 257988 7608
rect 258040 7596 258046 7608
rect 476942 7596 476948 7608
rect 258040 7568 476948 7596
rect 258040 7556 258046 7568
rect 476942 7556 476948 7568
rect 477000 7556 477006 7608
rect 248322 7488 248328 7540
rect 248380 7528 248386 7540
rect 437934 7528 437940 7540
rect 248380 7500 437940 7528
rect 248380 7488 248386 7500
rect 437934 7488 437940 7500
rect 437992 7488 437998 7540
rect 246942 7420 246948 7472
rect 247000 7460 247006 7472
rect 434438 7460 434444 7472
rect 247000 7432 434444 7460
rect 247000 7420 247006 7432
rect 434438 7420 434444 7432
rect 434496 7420 434502 7472
rect 245562 7352 245568 7404
rect 245620 7392 245626 7404
rect 430850 7392 430856 7404
rect 245620 7364 430856 7392
rect 245620 7352 245626 7364
rect 430850 7352 430856 7364
rect 430908 7352 430914 7404
rect 245470 7284 245476 7336
rect 245528 7324 245534 7336
rect 427262 7324 427268 7336
rect 245528 7296 427268 7324
rect 245528 7284 245534 7296
rect 427262 7284 427268 7296
rect 427320 7284 427326 7336
rect 244182 7216 244188 7268
rect 244240 7256 244246 7268
rect 423766 7256 423772 7268
rect 244240 7228 423772 7256
rect 244240 7216 244246 7228
rect 423766 7216 423772 7228
rect 423824 7216 423830 7268
rect 242710 7148 242716 7200
rect 242768 7188 242774 7200
rect 420178 7188 420184 7200
rect 242768 7160 420184 7188
rect 242768 7148 242774 7160
rect 420178 7148 420184 7160
rect 420236 7148 420242 7200
rect 242802 7080 242808 7132
rect 242860 7120 242866 7132
rect 416682 7120 416688 7132
rect 242860 7092 416688 7120
rect 242860 7080 242866 7092
rect 416682 7080 416688 7092
rect 416740 7080 416746 7132
rect 126974 7012 126980 7064
rect 127032 7052 127038 7064
rect 282914 7052 282920 7064
rect 127032 7024 282920 7052
rect 127032 7012 127038 7024
rect 282914 7012 282920 7024
rect 282972 7012 282978 7064
rect 283098 7012 283104 7064
rect 283156 7052 283162 7064
rect 323026 7052 323032 7064
rect 283156 7024 323032 7052
rect 283156 7012 283162 7024
rect 323026 7012 323032 7024
rect 323084 7012 323090 7064
rect 353110 7012 353116 7064
rect 353168 7052 353174 7064
rect 400122 7052 400128 7064
rect 353168 7024 400128 7052
rect 353168 7012 353174 7024
rect 400122 7012 400128 7024
rect 400180 7012 400186 7064
rect 261754 6808 261760 6860
rect 261812 6848 261818 6860
rect 298738 6848 298744 6860
rect 261812 6820 298744 6848
rect 261812 6808 261818 6820
rect 298738 6808 298744 6820
rect 298796 6808 298802 6860
rect 304350 6808 304356 6860
rect 304408 6848 304414 6860
rect 328454 6848 328460 6860
rect 304408 6820 328460 6848
rect 304408 6808 304414 6820
rect 328454 6808 328460 6820
rect 328512 6808 328518 6860
rect 347590 6808 347596 6860
rect 347648 6848 347654 6860
rect 378870 6848 378876 6860
rect 347648 6820 378876 6848
rect 347648 6808 347654 6820
rect 378870 6808 378876 6820
rect 378928 6808 378934 6860
rect 389818 6808 389824 6860
rect 389876 6848 389882 6860
rect 391842 6848 391848 6860
rect 389876 6820 391848 6848
rect 389876 6808 389882 6820
rect 391842 6808 391848 6820
rect 391900 6808 391906 6860
rect 519538 6808 519544 6860
rect 519596 6848 519602 6860
rect 580166 6848 580172 6860
rect 519596 6820 580172 6848
rect 519596 6808 519602 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 265342 6740 265348 6792
rect 265400 6780 265406 6792
rect 317506 6780 317512 6792
rect 265400 6752 317512 6780
rect 265400 6740 265406 6752
rect 317506 6740 317512 6752
rect 317564 6740 317570 6792
rect 318518 6740 318524 6792
rect 318576 6780 318582 6792
rect 331214 6780 331220 6792
rect 318576 6752 331220 6780
rect 318576 6740 318582 6752
rect 331214 6740 331220 6752
rect 331272 6740 331278 6792
rect 349062 6740 349068 6792
rect 349120 6780 349126 6792
rect 382366 6780 382372 6792
rect 349120 6752 382372 6780
rect 349120 6740 349126 6752
rect 382366 6740 382372 6752
rect 382424 6740 382430 6792
rect 390462 6740 390468 6792
rect 390520 6780 390526 6792
rect 545482 6780 545488 6792
rect 390520 6752 545488 6780
rect 390520 6740 390526 6752
rect 545482 6740 545488 6752
rect 545540 6740 545546 6792
rect 187326 6672 187332 6724
rect 187384 6712 187390 6724
rect 298094 6712 298100 6724
rect 187384 6684 298100 6712
rect 187384 6672 187390 6684
rect 298094 6672 298100 6684
rect 298152 6672 298158 6724
rect 300762 6672 300768 6724
rect 300820 6712 300826 6724
rect 327074 6712 327080 6724
rect 300820 6684 327080 6712
rect 300820 6672 300826 6684
rect 327074 6672 327080 6684
rect 327132 6672 327138 6724
rect 350350 6672 350356 6724
rect 350408 6712 350414 6724
rect 385954 6712 385960 6724
rect 350408 6684 385960 6712
rect 350408 6672 350414 6684
rect 385954 6672 385960 6684
rect 386012 6672 386018 6724
rect 391750 6672 391756 6724
rect 391808 6712 391814 6724
rect 549070 6712 549076 6724
rect 391808 6684 549076 6712
rect 391808 6672 391814 6684
rect 549070 6672 549076 6684
rect 549128 6672 549134 6724
rect 102226 6604 102232 6656
rect 102284 6644 102290 6656
rect 126238 6644 126244 6656
rect 102284 6616 126244 6644
rect 102284 6604 102290 6616
rect 126238 6604 126244 6616
rect 126296 6604 126302 6656
rect 166074 6604 166080 6656
rect 166132 6644 166138 6656
rect 287698 6644 287704 6656
rect 166132 6616 287704 6644
rect 166132 6604 166138 6616
rect 287698 6604 287704 6616
rect 287756 6604 287762 6656
rect 290182 6604 290188 6656
rect 290240 6644 290246 6656
rect 324314 6644 324320 6656
rect 290240 6616 324320 6644
rect 290240 6604 290246 6616
rect 324314 6604 324320 6616
rect 324372 6604 324378 6656
rect 350442 6604 350448 6656
rect 350500 6644 350506 6656
rect 389450 6644 389456 6656
rect 350500 6616 389456 6644
rect 350500 6604 350506 6616
rect 389450 6604 389456 6616
rect 389508 6604 389514 6656
rect 391658 6604 391664 6656
rect 391716 6644 391722 6656
rect 552658 6644 552664 6656
rect 391716 6616 552664 6644
rect 391716 6604 391722 6616
rect 552658 6604 552664 6616
rect 552716 6604 552722 6656
rect 98638 6536 98644 6588
rect 98696 6576 98702 6588
rect 125594 6576 125600 6588
rect 98696 6548 125600 6576
rect 98696 6536 98702 6548
rect 125594 6536 125600 6548
rect 125652 6536 125658 6588
rect 162486 6536 162492 6588
rect 162544 6576 162550 6588
rect 291194 6576 291200 6588
rect 162544 6548 291200 6576
rect 162544 6536 162550 6548
rect 291194 6536 291200 6548
rect 291252 6536 291258 6588
rect 293678 6536 293684 6588
rect 293736 6576 293742 6588
rect 325786 6576 325792 6588
rect 293736 6548 325792 6576
rect 293736 6536 293742 6548
rect 325786 6536 325792 6548
rect 325844 6536 325850 6588
rect 340782 6536 340788 6588
rect 340840 6576 340846 6588
rect 350350 6576 350356 6588
rect 340840 6548 350356 6576
rect 340840 6536 340846 6548
rect 350350 6536 350356 6548
rect 350408 6536 350414 6588
rect 351822 6536 351828 6588
rect 351880 6576 351886 6588
rect 393038 6576 393044 6588
rect 351880 6548 393044 6576
rect 351880 6536 351886 6548
rect 393038 6536 393044 6548
rect 393096 6536 393102 6588
rect 393222 6536 393228 6588
rect 393280 6576 393286 6588
rect 556154 6576 556160 6588
rect 393280 6548 556160 6576
rect 393280 6536 393286 6548
rect 556154 6536 556160 6548
rect 556212 6536 556218 6588
rect 95050 6468 95056 6520
rect 95108 6508 95114 6520
rect 124306 6508 124312 6520
rect 95108 6480 124312 6508
rect 95108 6468 95114 6480
rect 124306 6468 124312 6480
rect 124364 6468 124370 6520
rect 229002 6468 229008 6520
rect 229060 6508 229066 6520
rect 363506 6508 363512 6520
rect 229060 6480 363512 6508
rect 229060 6468 229066 6480
rect 363506 6468 363512 6480
rect 363564 6468 363570 6520
rect 394602 6468 394608 6520
rect 394660 6508 394666 6520
rect 559742 6508 559748 6520
rect 394660 6480 559748 6508
rect 394660 6468 394666 6480
rect 559742 6468 559748 6480
rect 559800 6468 559806 6520
rect 87966 6400 87972 6452
rect 88024 6440 88030 6452
rect 122834 6440 122840 6452
rect 88024 6412 122840 6440
rect 88024 6400 88030 6412
rect 122834 6400 122840 6412
rect 122892 6400 122898 6452
rect 230290 6400 230296 6452
rect 230348 6440 230354 6452
rect 367002 6440 367008 6452
rect 230348 6412 367008 6440
rect 230348 6400 230354 6412
rect 367002 6400 367008 6412
rect 367060 6400 367066 6452
rect 394510 6400 394516 6452
rect 394568 6440 394574 6452
rect 563238 6440 563244 6452
rect 394568 6412 563244 6440
rect 394568 6400 394574 6412
rect 563238 6400 563244 6412
rect 563296 6400 563302 6452
rect 63218 6332 63224 6384
rect 63276 6372 63282 6384
rect 116026 6372 116032 6384
rect 63276 6344 116032 6372
rect 63276 6332 63282 6344
rect 116026 6332 116032 6344
rect 116084 6332 116090 6384
rect 230382 6332 230388 6384
rect 230440 6372 230446 6384
rect 370590 6372 370596 6384
rect 230440 6344 370596 6372
rect 230440 6332 230446 6344
rect 370590 6332 370596 6344
rect 370648 6332 370654 6384
rect 371878 6332 371884 6384
rect 371936 6372 371942 6384
rect 384758 6372 384764 6384
rect 371936 6344 384764 6372
rect 371936 6332 371942 6344
rect 384758 6332 384764 6344
rect 384816 6332 384822 6384
rect 395982 6332 395988 6384
rect 396040 6372 396046 6384
rect 566826 6372 566832 6384
rect 396040 6344 566832 6372
rect 396040 6332 396046 6344
rect 566826 6332 566832 6344
rect 566884 6332 566890 6384
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 71038 6304 71044 6316
rect 2924 6276 71044 6304
rect 2924 6264 2930 6276
rect 71038 6264 71044 6276
rect 71096 6264 71102 6316
rect 71222 6264 71228 6316
rect 71280 6304 71286 6316
rect 146294 6304 146300 6316
rect 71280 6276 146300 6304
rect 71280 6264 71286 6276
rect 146294 6264 146300 6276
rect 146352 6264 146358 6316
rect 231670 6264 231676 6316
rect 231728 6304 231734 6316
rect 374086 6304 374092 6316
rect 231728 6276 374092 6304
rect 231728 6264 231734 6276
rect 374086 6264 374092 6276
rect 374144 6264 374150 6316
rect 392857 6307 392915 6313
rect 392857 6273 392869 6307
rect 392903 6304 392915 6307
rect 396534 6304 396540 6316
rect 392903 6276 396540 6304
rect 392903 6273 392915 6276
rect 392857 6267 392915 6273
rect 396534 6264 396540 6276
rect 396592 6264 396598 6316
rect 397270 6264 397276 6316
rect 397328 6304 397334 6316
rect 570322 6304 570328 6316
rect 397328 6276 570328 6304
rect 397328 6264 397334 6276
rect 570322 6264 570328 6276
rect 570380 6264 570386 6316
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 107654 6236 107660 6248
rect 27764 6208 107660 6236
rect 27764 6196 27770 6208
rect 107654 6196 107660 6208
rect 107712 6196 107718 6248
rect 116394 6196 116400 6248
rect 116452 6236 116458 6248
rect 129734 6236 129740 6248
rect 116452 6208 129740 6236
rect 116452 6196 116458 6208
rect 129734 6196 129740 6208
rect 129792 6196 129798 6248
rect 196618 6196 196624 6248
rect 196676 6236 196682 6248
rect 207382 6236 207388 6248
rect 196676 6208 207388 6236
rect 196676 6196 196682 6208
rect 207382 6196 207388 6208
rect 207440 6196 207446 6248
rect 231762 6196 231768 6248
rect 231820 6236 231826 6248
rect 377674 6236 377680 6248
rect 231820 6208 377680 6236
rect 231820 6196 231826 6208
rect 377674 6196 377680 6208
rect 377732 6196 377738 6248
rect 388990 6196 388996 6248
rect 389048 6236 389054 6248
rect 393961 6239 394019 6245
rect 393961 6236 393973 6239
rect 389048 6208 393973 6236
rect 389048 6196 389054 6208
rect 393961 6205 393973 6208
rect 394007 6205 394019 6239
rect 393961 6199 394019 6205
rect 397362 6196 397368 6248
rect 397420 6236 397426 6248
rect 573910 6236 573916 6248
rect 397420 6208 573916 6236
rect 397420 6196 397426 6208
rect 573910 6196 573916 6208
rect 573968 6196 573974 6248
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 106274 6168 106280 6180
rect 23072 6140 106280 6168
rect 23072 6128 23078 6140
rect 106274 6128 106280 6140
rect 106332 6128 106338 6180
rect 125870 6128 125876 6180
rect 125928 6168 125934 6180
rect 166258 6168 166264 6180
rect 125928 6140 166264 6168
rect 125928 6128 125934 6140
rect 166258 6128 166264 6140
rect 166316 6128 166322 6180
rect 186958 6128 186964 6180
rect 187016 6168 187022 6180
rect 196802 6168 196808 6180
rect 187016 6140 196808 6168
rect 187016 6128 187022 6140
rect 196802 6128 196808 6140
rect 196860 6128 196866 6180
rect 233142 6128 233148 6180
rect 233200 6168 233206 6180
rect 381170 6168 381176 6180
rect 233200 6140 381176 6168
rect 233200 6128 233206 6140
rect 381170 6128 381176 6140
rect 381228 6128 381234 6180
rect 387702 6128 387708 6180
rect 387760 6168 387766 6180
rect 390557 6171 390615 6177
rect 387760 6140 390508 6168
rect 387760 6128 387766 6140
rect 258718 6060 258724 6112
rect 258776 6100 258782 6112
rect 285398 6100 285404 6112
rect 258776 6072 285404 6100
rect 258776 6060 258782 6072
rect 285398 6060 285404 6072
rect 285456 6060 285462 6112
rect 286594 6060 286600 6112
rect 286652 6100 286658 6112
rect 322934 6100 322940 6112
rect 286652 6072 322940 6100
rect 286652 6060 286658 6072
rect 322934 6060 322940 6072
rect 322992 6060 322998 6112
rect 342070 6060 342076 6112
rect 342128 6100 342134 6112
rect 347593 6103 347651 6109
rect 347593 6100 347605 6103
rect 342128 6072 347605 6100
rect 342128 6060 342134 6072
rect 347593 6069 347605 6072
rect 347639 6069 347651 6103
rect 347593 6063 347651 6069
rect 347682 6060 347688 6112
rect 347740 6100 347746 6112
rect 375282 6100 375288 6112
rect 347740 6072 375288 6100
rect 347740 6060 347746 6072
rect 375282 6060 375288 6072
rect 375340 6060 375346 6112
rect 389082 6060 389088 6112
rect 389140 6100 389146 6112
rect 390373 6103 390431 6109
rect 390373 6100 390385 6103
rect 389140 6072 390385 6100
rect 389140 6060 389146 6072
rect 390373 6069 390385 6072
rect 390419 6069 390431 6103
rect 390373 6063 390431 6069
rect 264238 5992 264244 6044
rect 264296 6032 264302 6044
rect 292574 6032 292580 6044
rect 264296 6004 292580 6032
rect 264296 5992 264302 6004
rect 292574 5992 292580 6004
rect 292632 5992 292638 6044
rect 297266 5992 297272 6044
rect 297324 6032 297330 6044
rect 325694 6032 325700 6044
rect 297324 6004 325700 6032
rect 297324 5992 297330 6004
rect 325694 5992 325700 6004
rect 325752 5992 325758 6044
rect 346302 5992 346308 6044
rect 346360 6032 346366 6044
rect 371694 6032 371700 6044
rect 346360 6004 371700 6032
rect 346360 5992 346366 6004
rect 371694 5992 371700 6004
rect 371752 5992 371758 6044
rect 384942 5992 384948 6044
rect 385000 6032 385006 6044
rect 389177 6035 389235 6041
rect 389177 6032 389189 6035
rect 385000 6004 389189 6032
rect 385000 5992 385006 6004
rect 389177 6001 389189 6004
rect 389223 6001 389235 6035
rect 390480 6032 390508 6140
rect 390557 6137 390569 6171
rect 390603 6168 390615 6171
rect 390603 6140 394096 6168
rect 390603 6137 390615 6140
rect 390557 6131 390615 6137
rect 394068 6100 394096 6140
rect 398742 6128 398748 6180
rect 398800 6168 398806 6180
rect 577406 6168 577412 6180
rect 398800 6140 577412 6168
rect 398800 6128 398806 6140
rect 577406 6128 577412 6140
rect 577464 6128 577470 6180
rect 538398 6100 538404 6112
rect 394068 6072 538404 6100
rect 538398 6060 538404 6072
rect 538456 6060 538462 6112
rect 534902 6032 534908 6044
rect 390480 6004 534908 6032
rect 389177 5995 389235 6001
rect 534902 5992 534908 6004
rect 534960 5992 534966 6044
rect 284938 5924 284944 5976
rect 284996 5964 285002 5976
rect 299658 5964 299664 5976
rect 284996 5936 299664 5964
rect 284996 5924 285002 5936
rect 299658 5924 299664 5936
rect 299716 5924 299722 5976
rect 307938 5924 307944 5976
rect 307996 5964 308002 5976
rect 328546 5964 328552 5976
rect 307996 5936 328552 5964
rect 307996 5924 308002 5936
rect 328546 5924 328552 5936
rect 328604 5924 328610 5976
rect 344830 5924 344836 5976
rect 344888 5964 344894 5976
rect 368198 5964 368204 5976
rect 344888 5936 368204 5964
rect 344888 5924 344894 5936
rect 368198 5924 368204 5936
rect 368256 5924 368262 5976
rect 386230 5924 386236 5976
rect 386288 5964 386294 5976
rect 531314 5964 531320 5976
rect 386288 5936 531320 5964
rect 386288 5924 386294 5936
rect 531314 5924 531320 5936
rect 531372 5924 531378 5976
rect 311434 5856 311440 5908
rect 311492 5896 311498 5908
rect 329834 5896 329840 5908
rect 311492 5868 329840 5896
rect 311492 5856 311498 5868
rect 329834 5856 329840 5868
rect 329892 5856 329898 5908
rect 344922 5856 344928 5908
rect 344980 5896 344986 5908
rect 364610 5896 364616 5908
rect 344980 5868 364616 5896
rect 344980 5856 344986 5868
rect 364610 5856 364616 5868
rect 364668 5856 364674 5908
rect 386322 5856 386328 5908
rect 386380 5896 386386 5908
rect 527818 5896 527824 5908
rect 386380 5868 527824 5896
rect 386380 5856 386386 5868
rect 527818 5856 527824 5868
rect 527876 5856 527882 5908
rect 315022 5788 315028 5840
rect 315080 5828 315086 5840
rect 329926 5828 329932 5840
rect 315080 5800 329932 5828
rect 315080 5788 315086 5800
rect 329926 5788 329932 5800
rect 329984 5788 329990 5840
rect 343542 5788 343548 5840
rect 343600 5828 343606 5840
rect 361114 5828 361120 5840
rect 343600 5800 361120 5828
rect 343600 5788 343606 5800
rect 361114 5788 361120 5800
rect 361172 5788 361178 5840
rect 389177 5831 389235 5837
rect 389177 5797 389189 5831
rect 389223 5828 389235 5831
rect 524230 5828 524236 5840
rect 389223 5800 524236 5828
rect 389223 5797 389235 5800
rect 389177 5791 389235 5797
rect 524230 5788 524236 5800
rect 524288 5788 524294 5840
rect 322106 5720 322112 5772
rect 322164 5760 322170 5772
rect 332686 5760 332692 5772
rect 322164 5732 332692 5760
rect 322164 5720 322170 5732
rect 332686 5720 332692 5732
rect 332744 5720 332750 5772
rect 342162 5720 342168 5772
rect 342220 5760 342226 5772
rect 357526 5760 357532 5772
rect 342220 5732 357532 5760
rect 342220 5720 342226 5732
rect 357526 5720 357532 5732
rect 357584 5720 357590 5772
rect 383562 5720 383568 5772
rect 383620 5760 383626 5772
rect 520734 5760 520740 5772
rect 383620 5732 520740 5760
rect 383620 5720 383626 5732
rect 520734 5720 520740 5732
rect 520792 5720 520798 5772
rect 339402 5652 339408 5704
rect 339460 5692 339466 5704
rect 346946 5692 346952 5704
rect 339460 5664 346952 5692
rect 339460 5652 339466 5664
rect 346946 5652 346952 5664
rect 347004 5652 347010 5704
rect 347593 5695 347651 5701
rect 347593 5661 347605 5695
rect 347639 5692 347651 5695
rect 354030 5692 354036 5704
rect 347639 5664 354036 5692
rect 347639 5661 347651 5664
rect 347593 5655 347651 5661
rect 354030 5652 354036 5664
rect 354088 5652 354094 5704
rect 383470 5652 383476 5704
rect 383528 5692 383534 5704
rect 517146 5692 517152 5704
rect 383528 5664 517152 5692
rect 383528 5652 383534 5664
rect 517146 5652 517152 5664
rect 517204 5652 517210 5704
rect 332686 5584 332692 5636
rect 332744 5624 332750 5636
rect 335446 5624 335452 5636
rect 332744 5596 335452 5624
rect 332744 5584 332750 5596
rect 335446 5584 335452 5596
rect 335504 5584 335510 5636
rect 339310 5584 339316 5636
rect 339368 5624 339374 5636
rect 343358 5624 343364 5636
rect 339368 5596 343364 5624
rect 339368 5584 339374 5596
rect 343358 5584 343364 5596
rect 343416 5584 343422 5636
rect 382182 5584 382188 5636
rect 382240 5624 382246 5636
rect 513558 5624 513564 5636
rect 382240 5596 513564 5624
rect 382240 5584 382246 5596
rect 513558 5584 513564 5596
rect 513616 5584 513622 5636
rect 204898 5516 204904 5568
rect 204956 5556 204962 5568
rect 210970 5556 210976 5568
rect 204956 5528 210976 5556
rect 204956 5516 204962 5528
rect 210970 5516 210976 5528
rect 211028 5516 211034 5568
rect 329190 5516 329196 5568
rect 329248 5556 329254 5568
rect 333974 5556 333980 5568
rect 329248 5528 333980 5556
rect 329248 5516 329254 5528
rect 333974 5516 333980 5528
rect 334032 5516 334038 5568
rect 338022 5516 338028 5568
rect 338080 5556 338086 5568
rect 339862 5556 339868 5568
rect 338080 5528 339868 5556
rect 338080 5516 338086 5528
rect 339862 5516 339868 5528
rect 339920 5516 339926 5568
rect 353202 5516 353208 5568
rect 353260 5556 353266 5568
rect 392857 5559 392915 5565
rect 392857 5556 392869 5559
rect 353260 5528 392869 5556
rect 353260 5516 353266 5528
rect 392857 5525 392869 5528
rect 392903 5525 392915 5559
rect 392857 5519 392915 5525
rect 393961 5559 394019 5565
rect 393961 5525 393973 5559
rect 394007 5556 394019 5559
rect 541986 5556 541992 5568
rect 394007 5528 541992 5556
rect 394007 5525 394019 5528
rect 393961 5519 394019 5525
rect 541986 5516 541992 5528
rect 542044 5516 542050 5568
rect 100570 5448 100576 5500
rect 100628 5488 100634 5500
rect 111610 5488 111616 5500
rect 100628 5460 111616 5488
rect 100628 5448 100634 5460
rect 111610 5448 111616 5460
rect 111668 5448 111674 5500
rect 198550 5448 198556 5500
rect 198608 5488 198614 5500
rect 246298 5488 246304 5500
rect 198608 5460 246304 5488
rect 198608 5448 198614 5460
rect 246298 5448 246304 5460
rect 246356 5448 246362 5500
rect 274450 5448 274456 5500
rect 274508 5488 274514 5500
rect 540790 5488 540796 5500
rect 274508 5460 540796 5488
rect 274508 5448 274514 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 83274 5380 83280 5432
rect 83332 5420 83338 5432
rect 87598 5420 87604 5432
rect 83332 5392 87604 5420
rect 83332 5380 83338 5392
rect 87598 5380 87604 5392
rect 87656 5380 87662 5432
rect 102042 5380 102048 5432
rect 102100 5420 102106 5432
rect 115106 5420 115112 5432
rect 102100 5392 115112 5420
rect 102100 5380 102106 5392
rect 115106 5380 115112 5392
rect 115164 5380 115170 5432
rect 200022 5380 200028 5432
rect 200080 5420 200086 5432
rect 249978 5420 249984 5432
rect 200080 5392 249984 5420
rect 200080 5380 200086 5392
rect 249978 5380 249984 5392
rect 250036 5380 250042 5432
rect 274542 5380 274548 5432
rect 274600 5420 274606 5432
rect 544378 5420 544384 5432
rect 274600 5392 544384 5420
rect 274600 5380 274606 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 76190 5312 76196 5364
rect 76248 5352 76254 5364
rect 89806 5352 89812 5364
rect 76248 5324 89812 5352
rect 76248 5312 76254 5324
rect 89806 5312 89812 5324
rect 89864 5312 89870 5364
rect 105538 5312 105544 5364
rect 105596 5352 105602 5364
rect 122282 5352 122288 5364
rect 105596 5324 122288 5352
rect 105596 5312 105602 5324
rect 122282 5312 122288 5324
rect 122340 5312 122346 5364
rect 201402 5312 201408 5364
rect 201460 5352 201466 5364
rect 253474 5352 253480 5364
rect 201460 5324 253480 5352
rect 201460 5312 201466 5324
rect 253474 5312 253480 5324
rect 253532 5312 253538 5364
rect 254670 5312 254676 5364
rect 254728 5352 254734 5364
rect 262858 5352 262864 5364
rect 254728 5324 262864 5352
rect 254728 5312 254734 5324
rect 262858 5312 262864 5324
rect 262916 5312 262922 5364
rect 275922 5312 275928 5364
rect 275980 5352 275986 5364
rect 547874 5352 547880 5364
rect 275980 5324 547880 5352
rect 275980 5312 275986 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 72602 5244 72608 5296
rect 72660 5284 72666 5296
rect 86218 5284 86224 5296
rect 72660 5256 86224 5284
rect 72660 5244 72666 5256
rect 86218 5244 86224 5256
rect 86276 5244 86282 5296
rect 101950 5244 101956 5296
rect 102008 5284 102014 5296
rect 118786 5284 118792 5296
rect 102008 5256 118792 5284
rect 102008 5244 102014 5256
rect 118786 5244 118792 5256
rect 118844 5244 118850 5296
rect 201310 5244 201316 5296
rect 201368 5284 201374 5296
rect 257062 5284 257068 5296
rect 201368 5256 257068 5284
rect 201368 5244 201374 5256
rect 257062 5244 257068 5256
rect 257120 5244 257126 5296
rect 277302 5244 277308 5296
rect 277360 5284 277366 5296
rect 551462 5284 551468 5296
rect 277360 5256 551468 5284
rect 277360 5244 277366 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 59630 5176 59636 5228
rect 59688 5216 59694 5228
rect 79318 5216 79324 5228
rect 59688 5188 79324 5216
rect 59688 5176 59694 5188
rect 79318 5176 79324 5188
rect 79376 5176 79382 5228
rect 79686 5176 79692 5228
rect 79744 5216 79750 5228
rect 88978 5216 88984 5228
rect 79744 5188 88984 5216
rect 79744 5176 79750 5188
rect 88978 5176 88984 5188
rect 89036 5176 89042 5228
rect 91554 5176 91560 5228
rect 91612 5216 91618 5228
rect 123478 5216 123484 5228
rect 91612 5188 123484 5216
rect 91612 5176 91618 5188
rect 123478 5176 123484 5188
rect 123536 5176 123542 5228
rect 202782 5176 202788 5228
rect 202840 5216 202846 5228
rect 260650 5216 260656 5228
rect 202840 5188 260656 5216
rect 202840 5176 202846 5188
rect 260650 5176 260656 5188
rect 260708 5176 260714 5228
rect 277210 5176 277216 5228
rect 277268 5216 277274 5228
rect 554958 5216 554964 5228
rect 277268 5188 554964 5216
rect 277268 5176 277274 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 44266 5108 44272 5160
rect 44324 5148 44330 5160
rect 82814 5148 82820 5160
rect 44324 5120 82820 5148
rect 44324 5108 44330 5120
rect 82814 5108 82820 5120
rect 82872 5108 82878 5160
rect 84470 5108 84476 5160
rect 84528 5148 84534 5160
rect 121638 5148 121644 5160
rect 84528 5120 121644 5148
rect 84528 5108 84534 5120
rect 121638 5108 121644 5120
rect 121696 5108 121702 5160
rect 204162 5108 204168 5160
rect 204220 5148 204226 5160
rect 264146 5148 264152 5160
rect 204220 5120 264152 5148
rect 204220 5108 204226 5120
rect 264146 5108 264152 5120
rect 264204 5108 264210 5160
rect 279970 5108 279976 5160
rect 280028 5148 280034 5160
rect 282273 5151 282331 5157
rect 282273 5148 282285 5151
rect 280028 5120 282285 5148
rect 280028 5108 280034 5120
rect 282273 5117 282285 5120
rect 282319 5117 282331 5151
rect 282273 5111 282331 5117
rect 282365 5151 282423 5157
rect 282365 5117 282377 5151
rect 282411 5148 282423 5151
rect 558546 5148 558552 5160
rect 282411 5120 558552 5148
rect 282411 5117 282423 5120
rect 282365 5111 282423 5117
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 26510 5040 26516 5092
rect 26568 5080 26574 5092
rect 57238 5080 57244 5092
rect 26568 5052 57244 5080
rect 26568 5040 26574 5052
rect 57238 5040 57244 5052
rect 57296 5040 57302 5092
rect 66714 5040 66720 5092
rect 66772 5080 66778 5092
rect 116578 5080 116584 5092
rect 66772 5052 116584 5080
rect 66772 5040 66778 5052
rect 116578 5040 116584 5052
rect 116636 5040 116642 5092
rect 140038 5040 140044 5092
rect 140096 5080 140102 5092
rect 162118 5080 162124 5092
rect 140096 5052 162124 5080
rect 140096 5040 140102 5052
rect 162118 5040 162124 5052
rect 162176 5040 162182 5092
rect 204070 5040 204076 5092
rect 204128 5080 204134 5092
rect 267734 5080 267740 5092
rect 204128 5052 267740 5080
rect 204128 5040 204134 5052
rect 267734 5040 267740 5052
rect 267792 5040 267798 5092
rect 280062 5040 280068 5092
rect 280120 5080 280126 5092
rect 562042 5080 562048 5092
rect 280120 5052 562048 5080
rect 280120 5040 280126 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 34790 4972 34796 5024
rect 34848 5012 34854 5024
rect 50338 5012 50344 5024
rect 34848 4984 50344 5012
rect 34848 4972 34854 4984
rect 50338 4972 50344 4984
rect 50396 4972 50402 5024
rect 56042 4972 56048 5024
rect 56100 5012 56106 5024
rect 114646 5012 114652 5024
rect 56100 4984 114652 5012
rect 56100 4972 56106 4984
rect 114646 4972 114652 4984
rect 114704 4972 114710 5024
rect 147122 4972 147128 5024
rect 147180 5012 147186 5024
rect 172514 5012 172520 5024
rect 147180 4984 172520 5012
rect 147180 4972 147186 4984
rect 172514 4972 172520 4984
rect 172572 4972 172578 5024
rect 205542 4972 205548 5024
rect 205600 5012 205606 5024
rect 271230 5012 271236 5024
rect 205600 4984 271236 5012
rect 205600 4972 205606 4984
rect 271230 4972 271236 4984
rect 271288 4972 271294 5024
rect 271690 4972 271696 5024
rect 271748 5012 271754 5024
rect 282181 5015 282239 5021
rect 282181 5012 282193 5015
rect 271748 4984 282193 5012
rect 271748 4972 271754 4984
rect 282181 4981 282193 4984
rect 282227 4981 282239 5015
rect 282181 4975 282239 4981
rect 282273 5015 282331 5021
rect 282273 4981 282285 5015
rect 282319 5012 282331 5015
rect 565630 5012 565636 5024
rect 282319 4984 565636 5012
rect 282319 4981 282331 4984
rect 282273 4975 282331 4981
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 7650 4904 7656 4956
rect 7708 4944 7714 4956
rect 74626 4944 74632 4956
rect 7708 4916 74632 4944
rect 7708 4904 7714 4916
rect 74626 4904 74632 4916
rect 74684 4904 74690 4956
rect 77386 4904 77392 4956
rect 77444 4944 77450 4956
rect 115198 4944 115204 4956
rect 77444 4916 115204 4944
rect 77444 4904 77450 4916
rect 115198 4904 115204 4916
rect 115256 4904 115262 4956
rect 136542 4904 136548 4956
rect 136600 4944 136606 4956
rect 169754 4944 169760 4956
rect 136600 4916 169760 4944
rect 136600 4904 136606 4916
rect 169754 4904 169760 4916
rect 169812 4904 169818 4956
rect 184842 4904 184848 4956
rect 184900 4944 184906 4956
rect 193214 4944 193220 4956
rect 184900 4916 193220 4944
rect 184900 4904 184906 4916
rect 193214 4904 193220 4916
rect 193272 4904 193278 4956
rect 206830 4904 206836 4956
rect 206888 4944 206894 4956
rect 274818 4944 274824 4956
rect 206888 4916 274824 4944
rect 206888 4904 206894 4916
rect 274818 4904 274824 4916
rect 274876 4904 274882 4956
rect 281350 4904 281356 4956
rect 281408 4944 281414 4956
rect 569126 4944 569132 4956
rect 281408 4916 569132 4944
rect 281408 4904 281414 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 71866 4876 71872 4888
rect 624 4848 71872 4876
rect 624 4836 630 4848
rect 71866 4836 71872 4848
rect 71924 4836 71930 4888
rect 73798 4836 73804 4888
rect 73856 4876 73862 4888
rect 118878 4876 118884 4888
rect 73856 4848 118884 4876
rect 73856 4836 73862 4848
rect 118878 4836 118884 4848
rect 118936 4836 118942 4888
rect 123478 4836 123484 4888
rect 123536 4876 123542 4888
rect 132494 4876 132500 4888
rect 123536 4848 132500 4876
rect 123536 4836 123542 4848
rect 132494 4836 132500 4848
rect 132552 4836 132558 4888
rect 132954 4836 132960 4888
rect 133012 4876 133018 4888
rect 168374 4876 168380 4888
rect 133012 4848 168380 4876
rect 133012 4836 133018 4848
rect 168374 4836 168380 4848
rect 168432 4836 168438 4888
rect 191098 4836 191104 4888
rect 191156 4876 191162 4888
rect 200298 4876 200304 4888
rect 191156 4848 200304 4876
rect 191156 4836 191162 4848
rect 200298 4836 200304 4848
rect 200356 4836 200362 4888
rect 206922 4836 206928 4888
rect 206980 4876 206986 4888
rect 272521 4879 272579 4885
rect 272521 4876 272533 4879
rect 206980 4848 272533 4876
rect 206980 4836 206986 4848
rect 272521 4845 272533 4848
rect 272567 4845 272579 4879
rect 272521 4839 272579 4845
rect 272610 4836 272616 4888
rect 272668 4876 272674 4888
rect 278038 4876 278044 4888
rect 272668 4848 278044 4876
rect 272668 4836 272674 4848
rect 278038 4836 278044 4848
rect 278096 4836 278102 4888
rect 281442 4836 281448 4888
rect 281500 4876 281506 4888
rect 572714 4876 572720 4888
rect 281500 4848 572720 4876
rect 281500 4836 281506 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 103698 4808 103704 4820
rect 8812 4780 103704 4808
rect 8812 4768 8818 4780
rect 103698 4768 103704 4780
rect 103756 4768 103762 4820
rect 109310 4768 109316 4820
rect 109368 4808 109374 4820
rect 128354 4808 128360 4820
rect 109368 4780 128360 4808
rect 109368 4768 109374 4780
rect 128354 4768 128360 4780
rect 128412 4768 128418 4820
rect 129366 4768 129372 4820
rect 129424 4808 129430 4820
rect 168466 4808 168472 4820
rect 129424 4780 168472 4808
rect 129424 4768 129430 4780
rect 168466 4768 168472 4780
rect 168524 4768 168530 4820
rect 187602 4768 187608 4820
rect 187660 4808 187666 4820
rect 203886 4808 203892 4820
rect 187660 4780 203892 4808
rect 187660 4768 187666 4780
rect 203886 4768 203892 4780
rect 203944 4768 203950 4820
rect 208302 4768 208308 4820
rect 208360 4808 208366 4820
rect 281902 4808 281908 4820
rect 208360 4780 281908 4808
rect 208360 4768 208366 4780
rect 281902 4768 281908 4780
rect 281960 4768 281966 4820
rect 282822 4768 282828 4820
rect 282880 4808 282886 4820
rect 576302 4808 576308 4820
rect 282880 4780 576308 4808
rect 282880 4768 282886 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 99282 4700 99288 4752
rect 99340 4740 99346 4752
rect 108114 4740 108120 4752
rect 99340 4712 108120 4740
rect 99340 4700 99346 4712
rect 108114 4700 108120 4712
rect 108172 4700 108178 4752
rect 198642 4700 198648 4752
rect 198700 4740 198706 4752
rect 242894 4740 242900 4752
rect 198700 4712 242900 4740
rect 198700 4700 198706 4712
rect 242894 4700 242900 4712
rect 242952 4700 242958 4752
rect 272521 4743 272579 4749
rect 272521 4709 272533 4743
rect 272567 4740 272579 4743
rect 278314 4740 278320 4752
rect 272567 4712 278320 4740
rect 272567 4709 272579 4712
rect 272521 4703 272579 4709
rect 278314 4700 278320 4712
rect 278372 4700 278378 4752
rect 537202 4740 537208 4752
rect 278700 4712 537208 4740
rect 197262 4632 197268 4684
rect 197320 4672 197326 4684
rect 239306 4672 239312 4684
rect 197320 4644 239312 4672
rect 197320 4632 197326 4644
rect 239306 4632 239312 4644
rect 239364 4632 239370 4684
rect 273162 4632 273168 4684
rect 273220 4672 273226 4684
rect 278700 4672 278728 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 533706 4672 533712 4684
rect 273220 4644 278728 4672
rect 278792 4644 533712 4672
rect 273220 4632 273226 4644
rect 99190 4564 99196 4616
rect 99248 4604 99254 4616
rect 104526 4604 104532 4616
rect 99248 4576 104532 4604
rect 99248 4564 99254 4576
rect 104526 4564 104532 4576
rect 104584 4564 104590 4616
rect 195882 4564 195888 4616
rect 195940 4604 195946 4616
rect 235810 4604 235816 4616
rect 195940 4576 235816 4604
rect 195940 4564 195946 4576
rect 235810 4564 235816 4576
rect 235868 4564 235874 4616
rect 271782 4564 271788 4616
rect 271840 4604 271846 4616
rect 278792 4604 278820 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 271840 4576 278820 4604
rect 282181 4607 282239 4613
rect 271840 4564 271846 4576
rect 282181 4573 282193 4607
rect 282227 4604 282239 4607
rect 530118 4604 530124 4616
rect 282227 4576 530124 4604
rect 282227 4573 282239 4576
rect 282181 4567 282239 4573
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 90358 4496 90364 4548
rect 90416 4536 90422 4548
rect 93854 4536 93860 4548
rect 90416 4508 93860 4536
rect 90416 4496 90422 4508
rect 93854 4496 93860 4508
rect 93912 4496 93918 4548
rect 195790 4496 195796 4548
rect 195848 4536 195854 4548
rect 232222 4536 232228 4548
rect 195848 4508 232228 4536
rect 195848 4496 195854 4508
rect 232222 4496 232228 4508
rect 232280 4496 232286 4548
rect 270402 4496 270408 4548
rect 270460 4536 270466 4548
rect 526622 4536 526628 4548
rect 270460 4508 526628 4536
rect 270460 4496 270466 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 194502 4428 194508 4480
rect 194560 4468 194566 4480
rect 228726 4468 228732 4480
rect 194560 4440 228732 4468
rect 194560 4428 194566 4440
rect 228726 4428 228732 4440
rect 228784 4428 228790 4480
rect 268930 4428 268936 4480
rect 268988 4468 268994 4480
rect 523034 4468 523040 4480
rect 268988 4440 523040 4468
rect 268988 4428 268994 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 193122 4360 193128 4412
rect 193180 4400 193186 4412
rect 225138 4400 225144 4412
rect 193180 4372 225144 4400
rect 193180 4360 193186 4372
rect 225138 4360 225144 4372
rect 225196 4360 225202 4412
rect 269022 4360 269028 4412
rect 269080 4400 269086 4412
rect 519538 4400 519544 4412
rect 269080 4372 519544 4400
rect 269080 4360 269086 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 193030 4292 193036 4344
rect 193088 4332 193094 4344
rect 221550 4332 221556 4344
rect 193088 4304 221556 4332
rect 193088 4292 193094 4304
rect 221550 4292 221556 4304
rect 221608 4292 221614 4344
rect 267642 4292 267648 4344
rect 267700 4332 267706 4344
rect 515950 4332 515956 4344
rect 267700 4304 515956 4332
rect 267700 4292 267706 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 191742 4224 191748 4276
rect 191800 4264 191806 4276
rect 218054 4264 218060 4276
rect 191800 4236 218060 4264
rect 191800 4224 191806 4236
rect 218054 4224 218060 4236
rect 218112 4224 218118 4276
rect 266262 4224 266268 4276
rect 266320 4264 266326 4276
rect 512454 4264 512460 4276
rect 266320 4236 512460 4264
rect 266320 4224 266326 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 48958 4156 48964 4208
rect 49016 4196 49022 4208
rect 53098 4196 53104 4208
rect 49016 4168 53104 4196
rect 49016 4156 49022 4168
rect 53098 4156 53104 4168
rect 53156 4156 53162 4208
rect 86862 4156 86868 4208
rect 86920 4196 86926 4208
rect 92566 4196 92572 4208
rect 86920 4168 92572 4196
rect 86920 4156 86926 4168
rect 92566 4156 92572 4168
rect 92624 4156 92630 4208
rect 97902 4156 97908 4208
rect 97960 4196 97966 4208
rect 101030 4196 101036 4208
rect 97960 4168 101036 4196
rect 97960 4156 97966 4168
rect 101030 4156 101036 4168
rect 101088 4156 101094 4208
rect 188430 4156 188436 4208
rect 188488 4196 188494 4208
rect 189718 4196 189724 4208
rect 188488 4168 189724 4196
rect 188488 4156 188494 4168
rect 189718 4156 189724 4168
rect 189776 4156 189782 4208
rect 278682 4156 278688 4208
rect 278740 4196 278746 4208
rect 282365 4199 282423 4205
rect 282365 4196 282377 4199
rect 278740 4168 282377 4196
rect 278740 4156 278746 4168
rect 282365 4165 282377 4168
rect 282411 4165 282423 4199
rect 282365 4159 282423 4165
rect 407758 4156 407764 4208
rect 407816 4196 407822 4208
rect 409598 4196 409604 4208
rect 407816 4168 409604 4196
rect 407816 4156 407822 4168
rect 409598 4156 409604 4168
rect 409656 4156 409662 4208
rect 53742 4088 53748 4140
rect 53800 4128 53806 4140
rect 57330 4128 57336 4140
rect 53800 4100 57336 4128
rect 53800 4088 53806 4100
rect 57330 4088 57336 4100
rect 57388 4088 57394 4140
rect 64322 4088 64328 4140
rect 64380 4128 64386 4140
rect 65426 4128 65432 4140
rect 64380 4100 65432 4128
rect 64380 4088 64386 4100
rect 65426 4088 65432 4100
rect 65484 4088 65490 4140
rect 71498 4088 71504 4140
rect 71556 4128 71562 4140
rect 76558 4128 76564 4140
rect 71556 4100 76564 4128
rect 71556 4088 71562 4100
rect 76558 4088 76564 4100
rect 76616 4088 76622 4140
rect 89162 4088 89168 4140
rect 89220 4128 89226 4140
rect 89220 4100 151814 4128
rect 89220 4088 89226 4100
rect 45462 4020 45468 4072
rect 45520 4060 45526 4072
rect 51718 4060 51724 4072
rect 45520 4032 51724 4060
rect 45520 4020 45526 4032
rect 51718 4020 51724 4032
rect 51776 4020 51782 4072
rect 85666 4020 85672 4072
rect 85724 4060 85730 4072
rect 150434 4060 150440 4072
rect 85724 4032 150440 4060
rect 85724 4020 85730 4032
rect 150434 4020 150440 4032
rect 150492 4020 150498 4072
rect 151786 4004 151814 4100
rect 234614 4088 234620 4140
rect 234672 4128 234678 4140
rect 240870 4128 240876 4140
rect 234672 4100 240876 4128
rect 234672 4088 234678 4100
rect 240870 4088 240876 4100
rect 240928 4088 240934 4140
rect 344554 4088 344560 4140
rect 344612 4128 344618 4140
rect 377398 4128 377404 4140
rect 344612 4100 377404 4128
rect 344612 4088 344618 4100
rect 377398 4088 377404 4100
rect 377456 4088 377462 4140
rect 383562 4088 383568 4140
rect 383620 4128 383626 4140
rect 463878 4128 463884 4140
rect 383620 4100 463884 4128
rect 383620 4088 383626 4100
rect 463878 4088 463884 4100
rect 463936 4088 463942 4140
rect 489270 4088 489276 4140
rect 489328 4128 489334 4140
rect 491110 4128 491116 4140
rect 489328 4100 491116 4128
rect 489328 4088 489334 4100
rect 491110 4088 491116 4100
rect 491168 4088 491174 4140
rect 506290 4088 506296 4140
rect 506348 4128 506354 4140
rect 550266 4128 550272 4140
rect 506348 4100 550272 4128
rect 506348 4088 506354 4100
rect 550266 4088 550272 4100
rect 550324 4088 550330 4140
rect 255866 4020 255872 4072
rect 255924 4060 255930 4072
rect 269758 4060 269764 4072
rect 255924 4032 269764 4060
rect 255924 4020 255930 4032
rect 269758 4020 269764 4032
rect 269816 4020 269822 4072
rect 273622 4020 273628 4072
rect 273680 4060 273686 4072
rect 287790 4060 287796 4072
rect 273680 4032 287796 4060
rect 273680 4020 273686 4032
rect 287790 4020 287796 4032
rect 287848 4020 287854 4072
rect 340966 4020 340972 4072
rect 341024 4060 341030 4072
rect 376018 4060 376024 4072
rect 341024 4032 376024 4060
rect 341024 4020 341030 4032
rect 376018 4020 376024 4032
rect 376076 4020 376082 4072
rect 379974 4020 379980 4072
rect 380032 4060 380038 4072
rect 462314 4060 462320 4072
rect 380032 4032 462320 4060
rect 380032 4020 380038 4032
rect 462314 4020 462320 4032
rect 462372 4020 462378 4072
rect 507762 4020 507768 4072
rect 507820 4060 507826 4072
rect 553762 4060 553768 4072
rect 507820 4032 553768 4060
rect 507820 4020 507826 4032
rect 553762 4020 553768 4032
rect 553820 4020 553826 4072
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 18598 3992 18604 4004
rect 14792 3964 18604 3992
rect 14792 3952 14798 3964
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 50154 3952 50160 4004
rect 50212 3992 50218 4004
rect 58618 3992 58624 4004
rect 50212 3964 58624 3992
rect 50212 3952 50218 3964
rect 58618 3952 58624 3964
rect 58676 3952 58682 4004
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 150526 3992 150532 4004
rect 82136 3964 150532 3992
rect 82136 3952 82142 3964
rect 150526 3952 150532 3964
rect 150584 3952 150590 4004
rect 151786 3964 151820 4004
rect 151814 3952 151820 3964
rect 151872 3952 151878 4004
rect 151909 3995 151967 4001
rect 151909 3961 151921 3995
rect 151955 3992 151967 3995
rect 160370 3992 160376 4004
rect 151955 3964 160376 3992
rect 151955 3961 151967 3964
rect 151909 3955 151967 3961
rect 160370 3952 160376 3964
rect 160428 3952 160434 4004
rect 168374 3952 168380 4004
rect 168432 3992 168438 4004
rect 178034 3992 178040 4004
rect 168432 3964 178040 3992
rect 168432 3952 168438 3964
rect 178034 3952 178040 3964
rect 178092 3952 178098 4004
rect 216858 3952 216864 4004
rect 216916 3992 216922 4004
rect 220078 3992 220084 4004
rect 216916 3964 220084 3992
rect 216916 3952 216922 3964
rect 220078 3952 220084 3964
rect 220136 3952 220142 4004
rect 266538 3952 266544 4004
rect 266596 3992 266602 4004
rect 282178 3992 282184 4004
rect 266596 3964 282184 3992
rect 266596 3952 266602 3964
rect 282178 3952 282184 3964
rect 282236 3952 282242 4004
rect 305546 3952 305552 4004
rect 305604 3992 305610 4004
rect 316770 3992 316776 4004
rect 305604 3964 316776 3992
rect 305604 3952 305610 3964
rect 316770 3952 316776 3964
rect 316828 3952 316834 4004
rect 333882 3952 333888 4004
rect 333940 3992 333946 4004
rect 363598 3992 363604 4004
rect 333940 3964 363604 3992
rect 333940 3952 333946 3964
rect 363598 3952 363604 3964
rect 363656 3952 363662 4004
rect 376478 3952 376484 4004
rect 376536 3992 376542 4004
rect 461026 3992 461032 4004
rect 376536 3964 461032 3992
rect 376536 3952 376542 3964
rect 461026 3952 461032 3964
rect 461084 3952 461090 4004
rect 509050 3952 509056 4004
rect 509108 3992 509114 4004
rect 557350 3992 557356 4004
rect 509108 3964 557356 3992
rect 509108 3952 509114 3964
rect 557350 3952 557356 3964
rect 557408 3952 557414 4004
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 47578 3924 47584 3936
rect 38436 3896 47584 3924
rect 38436 3884 38442 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 57238 3884 57244 3936
rect 57296 3924 57302 3936
rect 68370 3924 68376 3936
rect 57296 3896 68376 3924
rect 57296 3884 57302 3896
rect 68370 3884 68376 3896
rect 68428 3884 68434 3936
rect 78582 3884 78588 3936
rect 78640 3924 78646 3936
rect 149054 3924 149060 3936
rect 78640 3896 149060 3924
rect 78640 3884 78646 3896
rect 149054 3884 149060 3896
rect 149112 3884 149118 3936
rect 157794 3884 157800 3936
rect 157852 3924 157858 3936
rect 175274 3924 175280 3936
rect 157852 3896 175280 3924
rect 157852 3884 157858 3896
rect 175274 3884 175280 3896
rect 175332 3884 175338 3936
rect 252370 3884 252376 3936
rect 252428 3924 252434 3936
rect 266998 3924 267004 3936
rect 252428 3896 267004 3924
rect 252428 3884 252434 3896
rect 266998 3884 267004 3896
rect 267056 3884 267062 3936
rect 277210 3884 277216 3936
rect 277268 3924 277274 3936
rect 291838 3924 291844 3936
rect 277268 3896 291844 3924
rect 277268 3884 277274 3896
rect 291838 3884 291844 3896
rect 291896 3884 291902 3936
rect 301958 3884 301964 3936
rect 302016 3924 302022 3936
rect 320818 3924 320824 3936
rect 302016 3896 320824 3924
rect 302016 3884 302022 3896
rect 320818 3884 320824 3896
rect 320876 3884 320882 3936
rect 330386 3884 330392 3936
rect 330444 3924 330450 3936
rect 360838 3924 360844 3936
rect 330444 3896 360844 3924
rect 330444 3884 330450 3896
rect 360838 3884 360844 3896
rect 360896 3884 360902 3936
rect 372890 3884 372896 3936
rect 372948 3924 372954 3936
rect 460934 3924 460940 3936
rect 372948 3896 460940 3924
rect 372948 3884 372954 3896
rect 460934 3884 460940 3896
rect 460992 3884 460998 3936
rect 509142 3884 509148 3936
rect 509200 3924 509206 3936
rect 560846 3924 560852 3936
rect 509200 3896 560852 3924
rect 509200 3884 509206 3896
rect 560846 3884 560852 3896
rect 560904 3884 560910 3936
rect 31294 3816 31300 3868
rect 31352 3856 31358 3868
rect 43438 3856 43444 3868
rect 31352 3828 43444 3856
rect 31352 3816 31358 3828
rect 43438 3816 43444 3828
rect 43496 3816 43502 3868
rect 46658 3816 46664 3868
rect 46716 3856 46722 3868
rect 140774 3856 140780 3868
rect 46716 3828 140780 3856
rect 46716 3816 46722 3828
rect 140774 3816 140780 3828
rect 140832 3816 140838 3868
rect 154206 3816 154212 3868
rect 154264 3856 154270 3868
rect 173894 3856 173900 3868
rect 154264 3828 173900 3856
rect 154264 3816 154270 3828
rect 173894 3816 173900 3828
rect 173952 3816 173958 3868
rect 227530 3816 227536 3868
rect 227588 3856 227594 3868
rect 238018 3856 238024 3868
rect 227588 3828 238024 3856
rect 227588 3816 227594 3828
rect 238018 3816 238024 3828
rect 238076 3816 238082 3868
rect 241698 3816 241704 3868
rect 241756 3856 241762 3868
rect 260098 3856 260104 3868
rect 241756 3828 260104 3856
rect 241756 3816 241762 3828
rect 260098 3816 260104 3828
rect 260156 3816 260162 3868
rect 270034 3816 270040 3868
rect 270092 3856 270098 3868
rect 289170 3856 289176 3868
rect 270092 3828 289176 3856
rect 270092 3816 270098 3828
rect 289170 3816 289176 3828
rect 289228 3816 289234 3868
rect 309042 3816 309048 3868
rect 309100 3856 309106 3868
rect 342898 3856 342904 3868
rect 309100 3828 342904 3856
rect 309100 3816 309106 3828
rect 342898 3816 342904 3828
rect 342956 3816 342962 3868
rect 369394 3816 369400 3868
rect 369452 3856 369458 3868
rect 451921 3859 451979 3865
rect 451921 3856 451933 3859
rect 369452 3828 451933 3856
rect 369452 3816 369458 3828
rect 451921 3825 451933 3828
rect 451967 3825 451979 3859
rect 458358 3856 458364 3868
rect 451921 3819 451979 3825
rect 452028 3828 458364 3856
rect 18230 3748 18236 3800
rect 18288 3788 18294 3800
rect 39298 3788 39304 3800
rect 18288 3760 39304 3788
rect 18288 3748 18294 3760
rect 39298 3748 39304 3760
rect 39356 3748 39362 3800
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 139394 3788 139400 3800
rect 43128 3760 139400 3788
rect 43128 3748 43134 3760
rect 139394 3748 139400 3760
rect 139452 3748 139458 3800
rect 150618 3748 150624 3800
rect 150676 3788 150682 3800
rect 173986 3788 173992 3800
rect 150676 3760 173992 3788
rect 150676 3748 150682 3760
rect 173986 3748 173992 3760
rect 174044 3748 174050 3800
rect 190822 3748 190828 3800
rect 190880 3788 190886 3800
rect 209038 3788 209044 3800
rect 190880 3760 209044 3788
rect 190880 3748 190886 3760
rect 209038 3748 209044 3760
rect 209096 3748 209102 3800
rect 238110 3748 238116 3800
rect 238168 3788 238174 3800
rect 249058 3788 249064 3800
rect 238168 3760 249064 3788
rect 238168 3748 238174 3760
rect 249058 3748 249064 3760
rect 249116 3748 249122 3800
rect 259454 3748 259460 3800
rect 259512 3788 259518 3800
rect 286318 3788 286324 3800
rect 259512 3760 286324 3788
rect 259512 3748 259518 3760
rect 286318 3748 286324 3760
rect 286376 3748 286382 3800
rect 294874 3748 294880 3800
rect 294932 3788 294938 3800
rect 318058 3788 318064 3800
rect 294932 3760 318064 3788
rect 294932 3748 294938 3760
rect 318058 3748 318064 3760
rect 318116 3748 318122 3800
rect 323302 3748 323308 3800
rect 323360 3788 323366 3800
rect 358170 3788 358176 3800
rect 323360 3760 358176 3788
rect 323360 3748 323366 3760
rect 358170 3748 358176 3760
rect 358228 3748 358234 3800
rect 365806 3748 365812 3800
rect 365864 3788 365870 3800
rect 452028 3788 452056 3828
rect 458358 3816 458364 3828
rect 458416 3816 458422 3868
rect 461305 3859 461363 3865
rect 461305 3825 461317 3859
rect 461351 3856 461363 3859
rect 472066 3856 472072 3868
rect 461351 3828 472072 3856
rect 461351 3825 461363 3828
rect 461305 3819 461363 3825
rect 472066 3816 472072 3828
rect 472124 3816 472130 3868
rect 495342 3816 495348 3868
rect 495400 3856 495406 3868
rect 504174 3856 504180 3868
rect 495400 3828 504180 3856
rect 495400 3816 495406 3828
rect 504174 3816 504180 3828
rect 504232 3816 504238 3868
rect 510522 3816 510528 3868
rect 510580 3856 510586 3868
rect 564434 3856 564440 3868
rect 510580 3828 564440 3856
rect 510580 3816 510586 3828
rect 564434 3816 564440 3828
rect 564492 3816 564498 3868
rect 365864 3760 452056 3788
rect 452120 3760 462268 3788
rect 365864 3748 365870 3760
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 134521 3723 134579 3729
rect 134521 3720 134533 3723
rect 39632 3692 134533 3720
rect 39632 3680 39638 3692
rect 134521 3689 134533 3692
rect 134567 3689 134579 3723
rect 134521 3683 134579 3689
rect 134613 3723 134671 3729
rect 134613 3689 134625 3723
rect 134659 3720 134671 3723
rect 136818 3720 136824 3732
rect 134659 3692 136824 3720
rect 134659 3689 134671 3692
rect 134613 3683 134671 3689
rect 136818 3680 136824 3692
rect 136876 3680 136882 3732
rect 160094 3680 160100 3732
rect 160152 3720 160158 3732
rect 405734 3720 405740 3732
rect 160152 3692 405740 3720
rect 160152 3680 160158 3692
rect 405734 3680 405740 3692
rect 405792 3680 405798 3732
rect 418982 3680 418988 3732
rect 419040 3720 419046 3732
rect 452120 3720 452148 3760
rect 419040 3692 452148 3720
rect 452197 3723 452255 3729
rect 419040 3680 419046 3692
rect 452197 3689 452209 3723
rect 452243 3720 452255 3723
rect 454405 3723 454463 3729
rect 454405 3720 454417 3723
rect 452243 3692 454417 3720
rect 452243 3689 452255 3692
rect 452197 3683 452255 3689
rect 454405 3689 454417 3692
rect 454451 3689 454463 3723
rect 454405 3683 454463 3689
rect 454494 3680 454500 3732
rect 454552 3720 454558 3732
rect 455322 3720 455328 3732
rect 454552 3692 455328 3720
rect 454552 3680 454558 3692
rect 455322 3680 455328 3692
rect 455380 3680 455386 3732
rect 455417 3723 455475 3729
rect 455417 3689 455429 3723
rect 455463 3720 455475 3723
rect 459554 3720 459560 3732
rect 455463 3692 459560 3720
rect 455463 3689 455475 3692
rect 455417 3683 455475 3689
rect 459554 3680 459560 3692
rect 459612 3680 459618 3732
rect 462240 3720 462268 3760
rect 468478 3748 468484 3800
rect 468536 3788 468542 3800
rect 495894 3788 495900 3800
rect 468536 3760 495900 3788
rect 468536 3748 468542 3760
rect 495894 3748 495900 3760
rect 495952 3748 495958 3800
rect 496630 3748 496636 3800
rect 496688 3788 496694 3800
rect 498381 3791 498439 3797
rect 498381 3788 498393 3791
rect 496688 3760 498393 3788
rect 496688 3748 496694 3760
rect 498381 3757 498393 3760
rect 498427 3757 498439 3791
rect 498381 3751 498439 3757
rect 511810 3748 511816 3800
rect 511868 3788 511874 3800
rect 568022 3788 568028 3800
rect 511868 3760 568028 3788
rect 511868 3748 511874 3760
rect 568022 3748 568028 3760
rect 568080 3748 568086 3800
rect 471974 3720 471980 3732
rect 462240 3692 471980 3720
rect 471974 3680 471980 3692
rect 472032 3680 472038 3732
rect 496722 3680 496728 3732
rect 496780 3720 496786 3732
rect 507670 3720 507676 3732
rect 496780 3692 507676 3720
rect 496780 3680 496786 3692
rect 507670 3680 507676 3692
rect 507728 3680 507734 3732
rect 511902 3680 511908 3732
rect 511960 3720 511966 3732
rect 571518 3720 571524 3732
rect 511960 3692 571524 3720
rect 511960 3680 511966 3692
rect 571518 3680 571524 3692
rect 571576 3680 571582 3732
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 35158 3652 35164 3664
rect 13596 3624 35164 3652
rect 13596 3612 13602 3624
rect 35158 3612 35164 3624
rect 35216 3612 35222 3664
rect 35986 3612 35992 3664
rect 36044 3652 36050 3664
rect 138014 3652 138020 3664
rect 36044 3624 138020 3652
rect 36044 3612 36050 3624
rect 138014 3612 138020 3624
rect 138072 3612 138078 3664
rect 156598 3612 156604 3664
rect 156656 3652 156662 3664
rect 405826 3652 405832 3664
rect 156656 3624 405832 3652
rect 156656 3612 156662 3624
rect 405826 3612 405832 3624
rect 405884 3612 405890 3664
rect 422570 3612 422576 3664
rect 422628 3652 422634 3664
rect 423582 3652 423588 3664
rect 422628 3624 423588 3652
rect 422628 3612 422634 3624
rect 423582 3612 423588 3624
rect 423640 3612 423646 3664
rect 429654 3612 429660 3664
rect 429712 3652 429718 3664
rect 430482 3652 430488 3664
rect 429712 3624 430488 3652
rect 429712 3612 429718 3624
rect 430482 3612 430488 3624
rect 430540 3612 430546 3664
rect 430577 3655 430635 3661
rect 430577 3621 430589 3655
rect 430623 3652 430635 3655
rect 461305 3655 461363 3661
rect 461305 3652 461317 3655
rect 430623 3624 461317 3652
rect 430623 3621 430635 3624
rect 430577 3615 430635 3621
rect 461305 3621 461317 3624
rect 461351 3621 461363 3655
rect 461305 3615 461363 3621
rect 461397 3655 461455 3661
rect 461397 3621 461409 3655
rect 461443 3652 461455 3655
rect 469306 3652 469312 3664
rect 461443 3624 469312 3652
rect 461443 3621 461455 3624
rect 461397 3615 461455 3621
rect 469306 3612 469312 3624
rect 469364 3612 469370 3664
rect 486418 3612 486424 3664
rect 486476 3652 486482 3664
rect 488810 3652 488816 3664
rect 486476 3624 488816 3652
rect 486476 3612 486482 3624
rect 488810 3612 488816 3624
rect 488868 3612 488874 3664
rect 489178 3612 489184 3664
rect 489236 3652 489242 3664
rect 494698 3652 494704 3664
rect 489236 3624 494704 3652
rect 489236 3612 489242 3624
rect 494698 3612 494704 3624
rect 494756 3612 494762 3664
rect 498102 3612 498108 3664
rect 498160 3652 498166 3664
rect 498381 3655 498439 3661
rect 498160 3624 498332 3652
rect 498160 3612 498166 3624
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 15838 3584 15844 3596
rect 10008 3556 15844 3584
rect 10008 3544 10014 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 29638 3584 29644 3596
rect 25372 3556 29644 3584
rect 25372 3544 25378 3556
rect 29638 3544 29644 3556
rect 29696 3544 29702 3596
rect 32490 3544 32496 3596
rect 32548 3584 32554 3596
rect 136634 3584 136640 3596
rect 32548 3556 136640 3584
rect 32548 3544 32554 3556
rect 136634 3544 136640 3556
rect 136692 3544 136698 3596
rect 151814 3544 151820 3596
rect 151872 3584 151878 3596
rect 153102 3584 153108 3596
rect 151872 3556 153108 3584
rect 151872 3544 151878 3556
rect 153102 3544 153108 3556
rect 153160 3544 153166 3596
rect 155402 3544 155408 3596
rect 155460 3584 155466 3596
rect 155862 3584 155868 3596
rect 155460 3556 155868 3584
rect 155460 3544 155466 3556
rect 155862 3544 155868 3556
rect 155920 3544 155926 3596
rect 158898 3544 158904 3596
rect 158956 3584 158962 3596
rect 160002 3584 160008 3596
rect 158956 3556 160008 3584
rect 158956 3544 158962 3556
rect 160002 3544 160008 3556
rect 160060 3544 160066 3596
rect 160097 3587 160155 3593
rect 160097 3553 160109 3587
rect 160143 3584 160155 3587
rect 404354 3584 404360 3596
rect 160143 3556 404360 3584
rect 160143 3553 160155 3556
rect 160097 3547 160155 3553
rect 404354 3544 404360 3556
rect 404412 3544 404418 3596
rect 411898 3544 411904 3596
rect 411956 3584 411962 3596
rect 470594 3584 470600 3596
rect 411956 3556 470600 3584
rect 411956 3544 411962 3556
rect 470594 3544 470600 3556
rect 470652 3544 470658 3596
rect 483750 3544 483756 3596
rect 483808 3584 483814 3596
rect 498194 3584 498200 3596
rect 483808 3556 498200 3584
rect 483808 3544 483814 3556
rect 498194 3544 498200 3556
rect 498252 3544 498258 3596
rect 498304 3584 498332 3624
rect 498381 3621 498393 3655
rect 498427 3652 498439 3655
rect 511258 3652 511264 3664
rect 498427 3624 511264 3652
rect 498427 3621 498439 3624
rect 498381 3615 498439 3621
rect 511258 3612 511264 3624
rect 511316 3612 511322 3664
rect 513282 3612 513288 3664
rect 513340 3652 513346 3664
rect 575106 3652 575112 3664
rect 513340 3624 575112 3652
rect 513340 3612 513346 3624
rect 575106 3612 575112 3624
rect 575164 3612 575170 3664
rect 514754 3584 514760 3596
rect 498304 3556 514760 3584
rect 514754 3544 514760 3556
rect 514812 3544 514818 3596
rect 517330 3544 517336 3596
rect 517388 3584 517394 3596
rect 582190 3584 582196 3596
rect 517388 3556 582196 3584
rect 517388 3544 517394 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4120 3488 16574 3516
rect 4120 3476 4126 3488
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 11698 3448 11704 3460
rect 1728 3420 11704 3448
rect 1728 3408 1734 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 16546 3448 16574 3488
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 25498 3516 25504 3528
rect 17972 3488 25504 3516
rect 17972 3448 18000 3488
rect 25498 3476 25504 3488
rect 25556 3476 25562 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 134613 3519 134671 3525
rect 134613 3516 134625 3519
rect 34624 3488 134625 3516
rect 16546 3420 18000 3448
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 24268 3420 26234 3448
rect 24268 3408 24274 3420
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 22738 3380 22744 3392
rect 15988 3352 22744 3380
rect 15988 3340 15994 3352
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 7558 3312 7564 3324
rect 6512 3284 7564 3312
rect 6512 3272 6518 3284
rect 7558 3272 7564 3284
rect 7616 3272 7622 3324
rect 26206 3312 26234 3420
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 34624 3380 34652 3488
rect 134613 3485 134625 3488
rect 134659 3485 134671 3519
rect 134613 3479 134671 3485
rect 134705 3519 134763 3525
rect 134705 3485 134717 3519
rect 134751 3516 134763 3519
rect 135165 3519 135223 3525
rect 135165 3516 135177 3519
rect 134751 3488 135177 3516
rect 134751 3485 134763 3488
rect 134705 3479 134763 3485
rect 135165 3485 135177 3488
rect 135211 3485 135223 3519
rect 135165 3479 135223 3485
rect 135254 3476 135260 3528
rect 135312 3516 135318 3528
rect 136450 3516 136456 3528
rect 135312 3488 136456 3516
rect 135312 3476 135318 3488
rect 136450 3476 136456 3488
rect 136508 3476 136514 3528
rect 138842 3476 138848 3528
rect 138900 3516 138906 3528
rect 139302 3516 139308 3528
rect 138900 3488 139308 3516
rect 138900 3476 138906 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 402974 3516 402980 3528
rect 149572 3488 402980 3516
rect 149572 3476 149578 3488
rect 402974 3476 402980 3488
rect 403032 3476 403038 3528
rect 408402 3476 408408 3528
rect 408460 3516 408466 3528
rect 408460 3488 461532 3516
rect 408460 3476 408466 3488
rect 135438 3448 135444 3460
rect 28960 3352 34652 3380
rect 35866 3420 135444 3448
rect 28960 3340 28966 3352
rect 35866 3312 35894 3420
rect 135438 3408 135444 3420
rect 135496 3408 135502 3460
rect 135533 3451 135591 3457
rect 135533 3417 135545 3451
rect 135579 3448 135591 3451
rect 139486 3448 139492 3460
rect 135579 3420 139492 3448
rect 135579 3417 135591 3420
rect 135533 3411 135591 3417
rect 139486 3408 139492 3420
rect 139544 3408 139550 3460
rect 142430 3408 142436 3460
rect 142488 3448 142494 3460
rect 143442 3448 143448 3460
rect 142488 3420 143448 3448
rect 142488 3408 142494 3420
rect 143442 3408 143448 3420
rect 143500 3408 143506 3460
rect 145926 3408 145932 3460
rect 145984 3448 145990 3460
rect 403066 3448 403072 3460
rect 145984 3420 403072 3448
rect 145984 3408 145990 3420
rect 403066 3408 403072 3420
rect 403124 3408 403130 3460
rect 404814 3408 404820 3460
rect 404872 3448 404878 3460
rect 461397 3451 461455 3457
rect 461397 3448 461409 3451
rect 404872 3420 461409 3448
rect 404872 3408 404878 3420
rect 461397 3417 461409 3420
rect 461443 3417 461455 3451
rect 461504 3448 461532 3488
rect 461578 3476 461584 3528
rect 461636 3516 461642 3528
rect 462222 3516 462228 3528
rect 461636 3488 462228 3516
rect 461636 3476 461642 3488
rect 462222 3476 462228 3488
rect 462280 3476 462286 3528
rect 465166 3476 465172 3528
rect 465224 3516 465230 3528
rect 466362 3516 466368 3528
rect 465224 3488 466368 3516
rect 465224 3476 465230 3488
rect 466362 3476 466368 3488
rect 466420 3476 466426 3528
rect 468662 3476 468668 3528
rect 468720 3516 468726 3528
rect 469122 3516 469128 3528
rect 468720 3488 469128 3516
rect 468720 3476 468726 3488
rect 469122 3476 469128 3488
rect 469180 3476 469186 3528
rect 472250 3476 472256 3528
rect 472308 3516 472314 3528
rect 473262 3516 473268 3528
rect 472308 3488 473268 3516
rect 472308 3476 472314 3488
rect 473262 3476 473268 3488
rect 473320 3476 473326 3528
rect 479334 3476 479340 3528
rect 479392 3516 479398 3528
rect 480162 3516 480168 3528
rect 479392 3488 480168 3516
rect 479392 3476 479398 3488
rect 480162 3476 480168 3488
rect 480220 3476 480226 3528
rect 486418 3476 486424 3528
rect 486476 3516 486482 3528
rect 487062 3516 487068 3528
rect 486476 3488 487068 3516
rect 486476 3476 486482 3488
rect 487062 3476 487068 3488
rect 487120 3476 487126 3528
rect 501598 3476 501604 3528
rect 501656 3516 501662 3528
rect 501656 3488 503116 3516
rect 501656 3476 501662 3488
rect 469398 3448 469404 3460
rect 461504 3420 469404 3448
rect 461397 3411 461455 3417
rect 469398 3408 469404 3420
rect 469456 3408 469462 3460
rect 471238 3408 471244 3460
rect 471296 3448 471302 3460
rect 502978 3448 502984 3460
rect 471296 3420 502984 3448
rect 471296 3408 471302 3420
rect 502978 3408 502984 3420
rect 503036 3408 503042 3460
rect 503088 3448 503116 3488
rect 504358 3476 504364 3528
rect 504416 3516 504422 3528
rect 505370 3516 505376 3528
rect 504416 3488 505376 3516
rect 504416 3476 504422 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 507118 3476 507124 3528
rect 507176 3516 507182 3528
rect 508866 3516 508872 3528
rect 507176 3488 508872 3516
rect 507176 3476 507182 3488
rect 508866 3476 508872 3488
rect 508924 3476 508930 3528
rect 514570 3476 514576 3528
rect 514628 3516 514634 3528
rect 578602 3516 578608 3528
rect 514628 3488 578608 3516
rect 514628 3476 514634 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 510062 3448 510068 3460
rect 503088 3420 510068 3448
rect 510062 3408 510068 3420
rect 510120 3408 510126 3460
rect 514662 3408 514668 3460
rect 514720 3448 514726 3460
rect 579798 3448 579804 3460
rect 514720 3420 579804 3448
rect 514720 3408 514726 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 42978 3380 42984 3392
rect 41932 3352 42984 3380
rect 41932 3340 41938 3352
rect 42978 3340 42984 3352
rect 43036 3340 43042 3392
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 52362 3380 52368 3392
rect 51408 3352 52368 3380
rect 51408 3340 51414 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 58434 3340 58440 3392
rect 58492 3380 58498 3392
rect 59262 3380 59268 3392
rect 58492 3352 59268 3380
rect 58492 3340 58498 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 60826 3340 60832 3392
rect 60884 3380 60890 3392
rect 61930 3380 61936 3392
rect 60884 3352 61936 3380
rect 60884 3340 60890 3352
rect 61930 3340 61936 3352
rect 61988 3340 61994 3392
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 66162 3380 66168 3392
rect 65576 3352 66168 3380
rect 65576 3340 65582 3352
rect 66162 3340 66168 3352
rect 66220 3340 66226 3392
rect 74994 3340 75000 3392
rect 75052 3380 75058 3392
rect 75822 3380 75828 3392
rect 75052 3352 75828 3380
rect 75052 3340 75058 3352
rect 75822 3340 75828 3352
rect 75880 3340 75886 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 92750 3340 92756 3392
rect 92808 3380 92814 3392
rect 92808 3352 152596 3380
rect 92808 3340 92814 3352
rect 26206 3284 35894 3312
rect 93946 3272 93952 3324
rect 94004 3312 94010 3324
rect 95142 3312 95148 3324
rect 94004 3284 95148 3312
rect 94004 3272 94010 3284
rect 95142 3272 95148 3284
rect 95200 3272 95206 3324
rect 99834 3272 99840 3324
rect 99892 3312 99898 3324
rect 100662 3312 100668 3324
rect 99892 3284 100668 3312
rect 99892 3272 99898 3284
rect 100662 3272 100668 3284
rect 100720 3272 100726 3324
rect 152568 3312 152596 3352
rect 153010 3340 153016 3392
rect 153068 3380 153074 3392
rect 160097 3383 160155 3389
rect 160097 3380 160109 3383
rect 153068 3352 160109 3380
rect 153068 3340 153074 3352
rect 160097 3349 160109 3352
rect 160143 3349 160155 3383
rect 160097 3343 160155 3349
rect 163682 3340 163688 3392
rect 163740 3380 163746 3392
rect 164142 3380 164148 3392
rect 163740 3352 164148 3380
rect 163740 3340 163746 3352
rect 164142 3340 164148 3352
rect 164200 3340 164206 3392
rect 164878 3340 164884 3392
rect 164936 3380 164942 3392
rect 165522 3380 165528 3392
rect 164936 3352 165528 3380
rect 164936 3340 164942 3352
rect 165522 3340 165528 3352
rect 165580 3340 165586 3392
rect 167178 3340 167184 3392
rect 167236 3380 167242 3392
rect 168282 3380 168288 3392
rect 167236 3352 168288 3380
rect 167236 3340 167242 3352
rect 168282 3340 168288 3352
rect 168340 3340 168346 3392
rect 173158 3340 173164 3392
rect 173216 3380 173222 3392
rect 173802 3380 173808 3392
rect 173216 3352 173808 3380
rect 173216 3340 173222 3352
rect 173802 3340 173808 3352
rect 173860 3340 173866 3392
rect 174262 3340 174268 3392
rect 174320 3380 174326 3392
rect 175182 3380 175188 3392
rect 174320 3352 175188 3380
rect 174320 3340 174326 3352
rect 175182 3340 175188 3352
rect 175240 3340 175246 3392
rect 180242 3340 180248 3392
rect 180300 3380 180306 3392
rect 180702 3380 180708 3392
rect 180300 3352 180708 3380
rect 180300 3340 180306 3352
rect 180702 3340 180708 3352
rect 180760 3340 180766 3392
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 182082 3380 182088 3392
rect 181496 3352 182088 3380
rect 181496 3340 181502 3352
rect 182082 3340 182088 3352
rect 182140 3340 182146 3392
rect 184934 3340 184940 3392
rect 184992 3380 184998 3392
rect 186222 3380 186228 3392
rect 184992 3352 186228 3380
rect 184992 3340 184998 3352
rect 186222 3340 186228 3352
rect 186280 3340 186286 3392
rect 188522 3340 188528 3392
rect 188580 3380 188586 3392
rect 188982 3380 188988 3392
rect 188580 3352 188988 3380
rect 188580 3340 188586 3352
rect 188982 3340 188988 3352
rect 189040 3340 189046 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 192938 3380 192944 3392
rect 192076 3352 192944 3380
rect 192076 3340 192082 3352
rect 192938 3340 192944 3352
rect 192996 3340 193002 3392
rect 199102 3340 199108 3392
rect 199160 3380 199166 3392
rect 199930 3380 199936 3392
rect 199160 3352 199936 3380
rect 199160 3340 199166 3352
rect 199930 3340 199936 3352
rect 199988 3340 199994 3392
rect 206186 3340 206192 3392
rect 206244 3380 206250 3392
rect 206738 3380 206744 3392
rect 206244 3352 206744 3380
rect 206244 3340 206250 3352
rect 206738 3340 206744 3352
rect 206796 3340 206802 3392
rect 209774 3340 209780 3392
rect 209832 3380 209838 3392
rect 211062 3380 211068 3392
rect 209832 3352 211068 3380
rect 209832 3340 209838 3352
rect 211062 3340 211068 3352
rect 211120 3340 211126 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 245194 3340 245200 3392
rect 245252 3380 245258 3392
rect 246390 3380 246396 3392
rect 245252 3352 246396 3380
rect 245252 3340 245258 3352
rect 246390 3340 246396 3352
rect 246448 3340 246454 3392
rect 258258 3340 258264 3392
rect 258316 3380 258322 3392
rect 259270 3380 259276 3392
rect 258316 3352 259276 3380
rect 258316 3340 258322 3352
rect 259270 3340 259276 3352
rect 259328 3340 259334 3392
rect 262950 3340 262956 3392
rect 263008 3380 263014 3392
rect 264330 3380 264336 3392
rect 263008 3352 264336 3380
rect 263008 3340 263014 3352
rect 264330 3340 264336 3352
rect 264388 3340 264394 3392
rect 276014 3340 276020 3392
rect 276072 3380 276078 3392
rect 277118 3380 277124 3392
rect 276072 3352 277124 3380
rect 276072 3340 276078 3352
rect 277118 3340 277124 3352
rect 277176 3340 277182 3392
rect 280706 3340 280712 3392
rect 280764 3380 280770 3392
rect 281258 3380 281264 3392
rect 280764 3352 281264 3380
rect 280764 3340 280770 3352
rect 281258 3340 281264 3352
rect 281316 3340 281322 3392
rect 291378 3340 291384 3392
rect 291436 3380 291442 3392
rect 292482 3380 292488 3392
rect 291436 3352 292488 3380
rect 291436 3340 291442 3352
rect 292482 3340 292488 3352
rect 292540 3340 292546 3392
rect 298462 3340 298468 3392
rect 298520 3380 298526 3392
rect 300118 3380 300124 3392
rect 298520 3352 300124 3380
rect 298520 3340 298526 3352
rect 300118 3340 300124 3352
rect 300176 3340 300182 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 319714 3340 319720 3392
rect 319772 3380 319778 3392
rect 323578 3380 323584 3392
rect 319772 3352 323584 3380
rect 319772 3340 319778 3352
rect 323578 3340 323584 3352
rect 323636 3340 323642 3392
rect 326798 3340 326804 3392
rect 326856 3380 326862 3392
rect 353938 3380 353944 3392
rect 326856 3352 353944 3380
rect 326856 3340 326862 3352
rect 353938 3340 353944 3352
rect 353996 3340 354002 3392
rect 387150 3340 387156 3392
rect 387208 3380 387214 3392
rect 463786 3380 463792 3392
rect 387208 3352 463792 3380
rect 387208 3340 387214 3352
rect 463786 3340 463792 3352
rect 463844 3340 463850 3392
rect 493962 3340 493968 3392
rect 494020 3380 494026 3392
rect 500586 3380 500592 3392
rect 494020 3352 500592 3380
rect 494020 3340 494026 3352
rect 500586 3340 500592 3352
rect 500644 3340 500650 3392
rect 506382 3340 506388 3392
rect 506440 3380 506446 3392
rect 546678 3380 546684 3392
rect 506440 3352 546684 3380
rect 506440 3340 506446 3352
rect 546678 3340 546684 3352
rect 546736 3340 546742 3392
rect 153286 3312 153292 3324
rect 100772 3284 152504 3312
rect 152568 3284 153292 3312
rect 96246 3204 96252 3256
rect 96304 3244 96310 3256
rect 100772 3244 100800 3284
rect 96304 3216 100800 3244
rect 96304 3204 96310 3216
rect 103330 3204 103336 3256
rect 103388 3244 103394 3256
rect 152476 3244 152504 3284
rect 153286 3272 153292 3284
rect 153344 3272 153350 3324
rect 175458 3272 175464 3324
rect 175516 3312 175522 3324
rect 179506 3312 179512 3324
rect 175516 3284 179512 3312
rect 175516 3272 175522 3284
rect 179506 3272 179512 3284
rect 179564 3272 179570 3324
rect 184198 3272 184204 3324
rect 184256 3312 184262 3324
rect 186130 3312 186136 3324
rect 184256 3284 186136 3312
rect 184256 3272 184262 3284
rect 186130 3272 186136 3284
rect 186188 3272 186194 3324
rect 287790 3272 287796 3324
rect 287848 3312 287854 3324
rect 294598 3312 294604 3324
rect 287848 3284 294604 3312
rect 287848 3272 287854 3284
rect 294598 3272 294604 3284
rect 294656 3272 294662 3324
rect 337470 3272 337476 3324
rect 337528 3312 337534 3324
rect 345658 3312 345664 3324
rect 337528 3284 345664 3312
rect 337528 3272 337534 3284
rect 345658 3272 345664 3284
rect 345716 3272 345722 3324
rect 348050 3272 348056 3324
rect 348108 3312 348114 3324
rect 374638 3312 374644 3324
rect 348108 3284 374644 3312
rect 348108 3272 348114 3284
rect 374638 3272 374644 3284
rect 374696 3272 374702 3324
rect 390646 3272 390652 3324
rect 390704 3312 390710 3324
rect 465258 3312 465264 3324
rect 390704 3284 465264 3312
rect 390704 3272 390710 3284
rect 465258 3272 465264 3284
rect 465316 3272 465322 3324
rect 505002 3272 505008 3324
rect 505060 3312 505066 3324
rect 543182 3312 543188 3324
rect 505060 3284 543188 3312
rect 505060 3272 505066 3284
rect 543182 3272 543188 3284
rect 543240 3272 543246 3324
rect 153194 3244 153200 3256
rect 103388 3216 152412 3244
rect 152476 3216 153200 3244
rect 103388 3204 103394 3216
rect 106918 3136 106924 3188
rect 106976 3176 106982 3188
rect 152384 3176 152412 3216
rect 153194 3204 153200 3216
rect 153252 3204 153258 3256
rect 171962 3204 171968 3256
rect 172020 3244 172026 3256
rect 177298 3244 177304 3256
rect 172020 3216 177304 3244
rect 172020 3204 172026 3216
rect 177298 3204 177304 3216
rect 177356 3204 177362 3256
rect 394234 3204 394240 3256
rect 394292 3244 394298 3256
rect 466638 3244 466644 3256
rect 394292 3216 466644 3244
rect 394292 3204 394298 3216
rect 466638 3204 466644 3216
rect 466696 3204 466702 3256
rect 503622 3204 503628 3256
rect 503680 3244 503686 3256
rect 539594 3244 539600 3256
rect 503680 3216 539600 3244
rect 503680 3204 503686 3216
rect 539594 3204 539600 3216
rect 539652 3204 539658 3256
rect 155954 3176 155960 3188
rect 106976 3148 152320 3176
rect 152384 3148 155960 3176
rect 106976 3136 106982 3148
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 14458 3108 14464 3120
rect 12400 3080 14464 3108
rect 12400 3068 12406 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 30098 3068 30104 3120
rect 30156 3108 30162 3120
rect 32398 3108 32404 3120
rect 30156 3080 32404 3108
rect 30156 3068 30162 3080
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 110506 3068 110512 3120
rect 110564 3108 110570 3120
rect 152292 3108 152320 3148
rect 155954 3136 155960 3148
rect 156012 3136 156018 3188
rect 183738 3136 183744 3188
rect 183796 3176 183802 3188
rect 188338 3176 188344 3188
rect 183796 3148 188344 3176
rect 183796 3136 183802 3148
rect 188338 3136 188344 3148
rect 188396 3136 188402 3188
rect 284294 3136 284300 3188
rect 284352 3176 284358 3188
rect 285582 3176 285588 3188
rect 284352 3148 285588 3176
rect 284352 3136 284358 3148
rect 285582 3136 285588 3148
rect 285640 3136 285646 3188
rect 316218 3136 316224 3188
rect 316276 3176 316282 3188
rect 322290 3176 322296 3188
rect 316276 3148 322296 3176
rect 316276 3136 316282 3148
rect 322290 3136 322296 3148
rect 322348 3136 322354 3188
rect 397730 3136 397736 3188
rect 397788 3176 397794 3188
rect 466546 3176 466552 3188
rect 397788 3148 466552 3176
rect 397788 3136 397794 3148
rect 466546 3136 466552 3148
rect 466604 3136 466610 3188
rect 493870 3136 493876 3188
rect 493928 3176 493934 3188
rect 497090 3176 497096 3188
rect 493928 3148 497096 3176
rect 493928 3136 493934 3148
rect 497090 3136 497096 3148
rect 497148 3136 497154 3188
rect 503530 3136 503536 3188
rect 503588 3176 503594 3188
rect 536098 3176 536104 3188
rect 503588 3148 536104 3176
rect 503588 3136 503594 3148
rect 536098 3136 536104 3148
rect 536156 3136 536162 3188
rect 156046 3108 156052 3120
rect 110564 3080 152228 3108
rect 152292 3080 156052 3108
rect 110564 3068 110570 3080
rect 67910 3000 67916 3052
rect 67968 3040 67974 3052
rect 71222 3040 71228 3052
rect 67968 3012 71228 3040
rect 67968 3000 67974 3012
rect 71222 3000 71228 3012
rect 71280 3000 71286 3052
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 152200 3040 152228 3080
rect 156046 3068 156052 3080
rect 156104 3068 156110 3120
rect 176654 3068 176660 3120
rect 176712 3108 176718 3120
rect 180058 3108 180064 3120
rect 176712 3080 180064 3108
rect 176712 3068 176718 3080
rect 180058 3068 180064 3080
rect 180116 3068 180122 3120
rect 231026 3068 231032 3120
rect 231084 3108 231090 3120
rect 233878 3108 233884 3120
rect 231084 3080 233884 3108
rect 231084 3068 231090 3080
rect 233878 3068 233884 3080
rect 233936 3068 233942 3120
rect 426158 3068 426164 3120
rect 426216 3108 426222 3120
rect 474826 3108 474832 3120
rect 426216 3080 474832 3108
rect 426216 3068 426222 3080
rect 474826 3068 474832 3080
rect 474884 3068 474890 3120
rect 485038 3068 485044 3120
rect 485096 3108 485102 3120
rect 487614 3108 487620 3120
rect 485096 3080 487620 3108
rect 485096 3068 485102 3080
rect 487614 3068 487620 3080
rect 487672 3068 487678 3120
rect 502242 3068 502248 3120
rect 502300 3108 502306 3120
rect 532510 3108 532516 3120
rect 502300 3080 532516 3108
rect 502300 3068 502306 3080
rect 532510 3068 532516 3080
rect 532568 3068 532574 3120
rect 157426 3040 157432 3052
rect 114060 3012 152136 3040
rect 152200 3012 157432 3040
rect 114060 3000 114066 3012
rect 117590 2932 117596 2984
rect 117648 2972 117654 2984
rect 152108 2972 152136 3012
rect 157426 3000 157432 3012
rect 157484 3000 157490 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 251818 3040 251824 3052
rect 248840 3012 251824 3040
rect 248840 3000 248846 3012
rect 251818 3000 251824 3012
rect 251876 3000 251882 3052
rect 415486 3000 415492 3052
rect 415544 3040 415550 3052
rect 430577 3043 430635 3049
rect 430577 3040 430589 3043
rect 415544 3012 430589 3040
rect 415544 3000 415550 3012
rect 430577 3009 430589 3012
rect 430623 3009 430635 3043
rect 476298 3040 476304 3052
rect 430577 3003 430635 3009
rect 441586 3012 476304 3040
rect 157334 2972 157340 2984
rect 117648 2944 152044 2972
rect 152108 2944 157340 2972
rect 117648 2932 117654 2944
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 151909 2907 151967 2913
rect 151909 2904 151921 2907
rect 121144 2876 151921 2904
rect 121144 2864 121150 2876
rect 151909 2873 151921 2876
rect 151955 2873 151967 2907
rect 152016 2904 152044 2944
rect 157334 2932 157340 2944
rect 157392 2932 157398 2984
rect 223942 2932 223948 2984
rect 224000 2972 224006 2984
rect 224770 2972 224776 2984
rect 224000 2944 224776 2972
rect 224000 2932 224006 2944
rect 224770 2932 224776 2944
rect 224828 2932 224834 2984
rect 433242 2932 433248 2984
rect 433300 2972 433306 2984
rect 441586 2972 441614 3012
rect 476298 3000 476304 3012
rect 476356 3000 476362 3052
rect 497458 3000 497464 3052
rect 497516 3040 497522 3052
rect 499390 3040 499396 3052
rect 497516 3012 499396 3040
rect 497516 3000 497522 3012
rect 499390 3000 499396 3012
rect 499448 3000 499454 3052
rect 500862 3000 500868 3052
rect 500920 3040 500926 3052
rect 529014 3040 529020 3052
rect 500920 3012 529020 3040
rect 500920 3000 500926 3012
rect 529014 3000 529020 3012
rect 529072 3000 529078 3052
rect 433300 2944 441614 2972
rect 433300 2932 433306 2944
rect 447410 2932 447416 2984
rect 447468 2972 447474 2984
rect 448422 2972 448428 2984
rect 447468 2944 448428 2972
rect 447468 2932 447474 2944
rect 448422 2932 448428 2944
rect 448480 2932 448486 2984
rect 476206 2972 476212 2984
rect 448532 2944 476212 2972
rect 158806 2904 158812 2916
rect 152016 2876 158812 2904
rect 151909 2867 151967 2873
rect 158806 2864 158812 2876
rect 158864 2864 158870 2916
rect 436738 2864 436744 2916
rect 436796 2904 436802 2916
rect 448532 2904 448560 2944
rect 476206 2932 476212 2944
rect 476264 2932 476270 2984
rect 490558 2932 490564 2984
rect 490616 2972 490622 2984
rect 492306 2972 492312 2984
rect 490616 2944 492312 2972
rect 490616 2932 490622 2944
rect 492306 2932 492312 2944
rect 492364 2932 492370 2984
rect 500770 2932 500776 2984
rect 500828 2972 500834 2984
rect 525426 2972 525432 2984
rect 500828 2944 525432 2972
rect 500828 2932 500834 2944
rect 525426 2932 525432 2944
rect 525484 2932 525490 2984
rect 478966 2904 478972 2916
rect 436796 2876 448560 2904
rect 448624 2876 478972 2904
rect 436796 2864 436802 2876
rect 124674 2796 124680 2848
rect 124732 2836 124738 2848
rect 160186 2836 160192 2848
rect 124732 2808 160192 2836
rect 124732 2796 124738 2808
rect 160186 2796 160192 2808
rect 160244 2796 160250 2848
rect 440326 2796 440332 2848
rect 440384 2836 440390 2848
rect 441522 2836 441528 2848
rect 440384 2808 441528 2836
rect 440384 2796 440390 2808
rect 441522 2796 441528 2808
rect 441580 2796 441586 2848
rect 443822 2796 443828 2848
rect 443880 2836 443886 2848
rect 448624 2836 448652 2876
rect 478966 2864 478972 2876
rect 479024 2864 479030 2916
rect 499482 2864 499488 2916
rect 499540 2904 499546 2916
rect 521838 2904 521844 2916
rect 499540 2876 521844 2904
rect 499540 2864 499546 2876
rect 521838 2864 521844 2876
rect 521896 2864 521902 2916
rect 443880 2808 448652 2836
rect 443880 2796 443886 2808
rect 450906 2796 450912 2848
rect 450964 2836 450970 2848
rect 480254 2836 480260 2848
rect 450964 2808 480260 2836
rect 450964 2796 450970 2808
rect 480254 2796 480260 2808
rect 480312 2796 480318 2848
rect 499298 2796 499304 2848
rect 499356 2836 499362 2848
rect 518342 2836 518348 2848
rect 499356 2808 518348 2836
rect 499356 2796 499362 2808
rect 518342 2796 518348 2808
rect 518400 2796 518406 2848
rect 340874 1912 340880 1964
rect 340932 1952 340938 1964
rect 342162 1952 342168 1964
rect 340932 1924 342168 1952
rect 340932 1912 340938 1924
rect 342162 1912 342168 1924
rect 342220 1912 342226 1964
<< via1 >>
rect 480168 700476 480220 700528
rect 527180 700476 527232 700528
rect 402888 700408 402940 700460
rect 429844 700408 429896 700460
rect 441528 700408 441580 700460
rect 478512 700408 478564 700460
rect 492588 700408 492640 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 378048 700340 378100 700392
rect 397460 700340 397512 700392
rect 416688 700340 416740 700392
rect 446128 700340 446180 700392
rect 453948 700340 454000 700392
rect 494796 700340 494848 700392
rect 505008 700340 505060 700392
rect 559656 700340 559708 700392
rect 339408 700272 339460 700324
rect 348792 700272 348844 700324
rect 351828 700272 351880 700324
rect 364984 700272 365036 700324
rect 365628 700272 365680 700324
rect 381176 700272 381228 700324
rect 390468 700272 390520 700324
rect 413652 700272 413704 700324
rect 429108 700272 429160 700324
rect 462320 700272 462372 700324
rect 466368 700272 466420 700324
rect 510988 700272 511040 700324
rect 517428 700272 517480 700324
rect 575848 700272 575900 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 56784 700136 56836 700188
rect 57888 700136 57940 700188
rect 186504 700136 186556 700188
rect 187608 700136 187660 700188
rect 251456 700068 251508 700120
rect 252468 700068 252520 700120
rect 283840 700068 283892 700120
rect 284944 700068 284996 700120
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 314568 699660 314620 699712
rect 316316 699660 316368 699712
rect 327724 699660 327776 699712
rect 332508 699660 332560 699712
rect 519544 696940 519596 696992
rect 580172 696940 580224 696992
rect 519636 683136 519688 683188
rect 580172 683136 580224 683188
rect 519728 670692 519780 670744
rect 580172 670692 580224 670744
rect 519820 656888 519872 656940
rect 580172 656888 580224 656940
rect 519912 643084 519964 643136
rect 580172 643084 580224 643136
rect 284944 643016 284996 643068
rect 288164 643016 288216 643068
rect 57888 642540 57940 642592
rect 110144 642540 110196 642592
rect 122748 642540 122800 642592
rect 161020 642540 161072 642592
rect 440884 642540 440936 642592
rect 441528 642540 441580 642592
rect 41328 642472 41380 642524
rect 97356 642472 97408 642524
rect 106188 642472 106240 642524
rect 148232 642472 148284 642524
rect 171048 642472 171100 642524
rect 199108 642472 199160 642524
rect 24768 642404 24820 642456
rect 84660 642404 84712 642456
rect 89628 642404 89680 642456
rect 135536 642404 135588 642456
rect 154488 642404 154540 642456
rect 186412 642404 186464 642456
rect 202788 642404 202840 642456
rect 224592 642404 224644 642456
rect 235908 642404 235960 642456
rect 249984 642404 250036 642456
rect 8208 642336 8260 642388
rect 72792 642336 72844 642388
rect 73068 642336 73120 642388
rect 122840 642336 122892 642388
rect 137928 642336 137980 642388
rect 173716 642336 173768 642388
rect 187608 642336 187660 642388
rect 211896 642336 211948 642388
rect 219348 642336 219400 642388
rect 237288 642336 237340 642388
rect 252468 642336 252520 642388
rect 262772 642336 262824 642388
rect 267648 642336 267700 642388
rect 275468 642336 275520 642388
rect 313648 641724 313700 641776
rect 314568 641724 314620 641776
rect 326344 641724 326396 641776
rect 327724 641724 327776 641776
rect 364524 641724 364576 641776
rect 365628 641724 365680 641776
rect 377220 641724 377272 641776
rect 378048 641724 378100 641776
rect 390008 641724 390060 641776
rect 390468 641724 390520 641776
rect 415400 641724 415452 641776
rect 416688 641724 416740 641776
rect 428096 641724 428148 641776
rect 429108 641724 429160 641776
rect 478972 641724 479024 641776
rect 480168 641724 480220 641776
rect 491760 641724 491812 641776
rect 492588 641724 492640 641776
rect 504456 641724 504508 641776
rect 505008 641724 505060 641776
rect 516508 641724 516560 641776
rect 517428 641724 517480 641776
rect 3424 637508 3476 637560
rect 69020 637508 69072 637560
rect 519544 630640 519596 630692
rect 580172 630640 580224 630692
rect 3516 626492 3568 626544
rect 69020 626492 69072 626544
rect 519636 616836 519688 616888
rect 580172 616836 580224 616888
rect 3608 615408 3660 615460
rect 69020 615408 69072 615460
rect 3700 605752 3752 605804
rect 69020 605752 69072 605804
rect 519728 603100 519780 603152
rect 580172 603100 580224 603152
rect 3792 594736 3844 594788
rect 69020 594736 69072 594788
rect 519820 590656 519872 590708
rect 579804 590656 579856 590708
rect 3424 583652 3476 583704
rect 69020 583652 69072 583704
rect 519544 576852 519596 576904
rect 580172 576852 580224 576904
rect 3516 572636 3568 572688
rect 69020 572636 69072 572688
rect 519636 563048 519688 563100
rect 579804 563048 579856 563100
rect 3608 561620 3660 561672
rect 69020 561620 69072 561672
rect 519728 550604 519780 550656
rect 580172 550604 580224 550656
rect 3700 550536 3752 550588
rect 69020 550536 69072 550588
rect 3424 539520 3476 539572
rect 69020 539520 69072 539572
rect 519820 536800 519872 536852
rect 580172 536800 580224 536852
rect 3516 528504 3568 528556
rect 69020 528504 69072 528556
rect 519544 524424 519596 524476
rect 580172 524424 580224 524476
rect 3608 517420 3660 517472
rect 69020 517420 69072 517472
rect 519636 510620 519688 510672
rect 580172 510620 580224 510672
rect 3700 507764 3752 507816
rect 69020 507764 69072 507816
rect 519728 496816 519780 496868
rect 580172 496816 580224 496868
rect 3424 496748 3476 496800
rect 69020 496748 69072 496800
rect 3516 485732 3568 485784
rect 69020 485732 69072 485784
rect 519544 484372 519596 484424
rect 580172 484372 580224 484424
rect 3608 474648 3660 474700
rect 69020 474648 69072 474700
rect 519636 470568 519688 470620
rect 579988 470568 580040 470620
rect 3424 463632 3476 463684
rect 69020 463632 69072 463684
rect 519544 456764 519596 456816
rect 580172 456764 580224 456816
rect 3516 452548 3568 452600
rect 69020 452548 69072 452600
rect 519636 444388 519688 444440
rect 580172 444388 580224 444440
rect 3608 441532 3660 441584
rect 69020 441532 69072 441584
rect 519544 430584 519596 430636
rect 580172 430584 580224 430636
rect 3424 430516 3476 430568
rect 69020 430516 69072 430568
rect 3516 419432 3568 419484
rect 69020 419432 69072 419484
rect 519636 418140 519688 418192
rect 580172 418140 580224 418192
rect 3424 409776 3476 409828
rect 69020 409776 69072 409828
rect 519544 404336 519596 404388
rect 580172 404336 580224 404388
rect 3516 398760 3568 398812
rect 69020 398760 69072 398812
rect 519544 390532 519596 390584
rect 580172 390532 580224 390584
rect 3424 387744 3476 387796
rect 69020 387744 69072 387796
rect 519544 378156 519596 378208
rect 580172 378156 580224 378208
rect 3424 376660 3476 376712
rect 69020 376660 69072 376712
rect 3424 365644 3476 365696
rect 69020 365644 69072 365696
rect 519360 364352 519412 364404
rect 580172 364352 580224 364404
rect 3424 354628 3476 354680
rect 69020 354628 69072 354680
rect 519820 351908 519872 351960
rect 580172 351908 580224 351960
rect 3148 343544 3200 343596
rect 69020 343544 69072 343596
rect 520004 338104 520056 338156
rect 580172 338104 580224 338156
rect 3424 331848 3476 331900
rect 69020 331848 69072 331900
rect 519360 325592 519412 325644
rect 580172 325592 580224 325644
rect 3424 320152 3476 320204
rect 69020 320152 69072 320204
rect 520188 313216 520240 313268
rect 580172 313216 580224 313268
rect 3424 309136 3476 309188
rect 69020 309136 69072 309188
rect 3424 299480 3476 299532
rect 69020 299480 69072 299532
rect 519360 299412 519412 299464
rect 580172 299412 580224 299464
rect 3424 288396 3476 288448
rect 69020 288396 69072 288448
rect 519544 285608 519596 285660
rect 580172 285608 580224 285660
rect 3516 277380 3568 277432
rect 69020 277380 69072 277432
rect 519544 273164 519596 273216
rect 580172 273164 580224 273216
rect 3424 266364 3476 266416
rect 69020 266364 69072 266416
rect 519544 259360 519596 259412
rect 580172 259360 580224 259412
rect 3516 255280 3568 255332
rect 69020 255280 69072 255332
rect 519636 245556 519688 245608
rect 580172 245556 580224 245608
rect 3424 244264 3476 244316
rect 69020 244264 69072 244316
rect 3516 233248 3568 233300
rect 69020 233248 69072 233300
rect 519544 233180 519596 233232
rect 579988 233180 580040 233232
rect 3424 222164 3476 222216
rect 69020 222164 69072 222216
rect 519636 219376 519688 219428
rect 580172 219376 580224 219428
rect 3608 211148 3660 211200
rect 69020 211148 69072 211200
rect 519544 206932 519596 206984
rect 579804 206932 579856 206984
rect 3516 201492 3568 201544
rect 69020 201492 69072 201544
rect 519728 193128 519780 193180
rect 580172 193128 580224 193180
rect 3424 190476 3476 190528
rect 69020 190476 69072 190528
rect 3608 179392 3660 179444
rect 69020 179392 69072 179444
rect 519636 179324 519688 179376
rect 580172 179324 580224 179376
rect 3516 168376 3568 168428
rect 69020 168376 69072 168428
rect 519544 166948 519596 167000
rect 580172 166948 580224 167000
rect 3424 157360 3476 157412
rect 69020 157360 69072 157412
rect 519728 153144 519780 153196
rect 580172 153144 580224 153196
rect 3700 146276 3752 146328
rect 69020 146276 69072 146328
rect 519636 139340 519688 139392
rect 580172 139340 580224 139392
rect 3608 135260 3660 135312
rect 69020 135260 69072 135312
rect 519544 126896 519596 126948
rect 580172 126896 580224 126948
rect 3516 124176 3568 124228
rect 69020 124176 69072 124228
rect 3424 113160 3476 113212
rect 69020 113160 69072 113212
rect 519820 113092 519872 113144
rect 579804 113092 579856 113144
rect 3792 103504 3844 103556
rect 69020 103504 69072 103556
rect 519728 100648 519780 100700
rect 580172 100648 580224 100700
rect 3700 92488 3752 92540
rect 69020 92488 69072 92540
rect 519636 86912 519688 86964
rect 580172 86912 580224 86964
rect 3608 81404 3660 81456
rect 69020 81404 69072 81456
rect 519544 73108 519596 73160
rect 580172 73108 580224 73160
rect 3516 70388 3568 70440
rect 69020 70388 69072 70440
rect 519912 60664 519964 60716
rect 580172 60664 580224 60716
rect 303620 59848 303672 59900
rect 304934 59848 304986 59900
rect 86960 59780 87012 59832
rect 88214 59780 88266 59832
rect 89812 59780 89864 59832
rect 90934 59780 90986 59832
rect 110420 59780 110472 59832
rect 111694 59780 111746 59832
rect 133972 59780 134024 59832
rect 135174 59780 135226 59832
rect 136640 59780 136692 59832
rect 137874 59780 137926 59832
rect 139400 59780 139452 59832
rect 140594 59780 140646 59832
rect 142160 59780 142212 59832
rect 143294 59780 143346 59832
rect 150440 59780 150492 59832
rect 151434 59780 151486 59832
rect 157340 59780 157392 59832
rect 158654 59780 158706 59832
rect 160192 59780 160244 59832
rect 161354 59780 161406 59832
rect 162952 59780 163004 59832
rect 164074 59780 164126 59832
rect 168380 59780 168432 59832
rect 169494 59780 169546 59832
rect 173900 59780 173952 59832
rect 174914 59780 174966 59832
rect 291200 59780 291252 59832
rect 292294 59780 292346 59832
rect 402980 59780 403032 59832
rect 404274 59780 404326 59832
rect 405740 59780 405792 59832
rect 406974 59780 407026 59832
rect 411260 59780 411312 59832
rect 412394 59780 412446 59832
rect 414020 59780 414072 59832
rect 415114 59780 415166 59832
rect 416780 59780 416832 59832
rect 417814 59780 417866 59832
rect 419540 59780 419592 59832
rect 420514 59780 420566 59832
rect 429200 59780 429252 59832
rect 430454 59780 430506 59832
rect 431960 59780 432012 59832
rect 433174 59780 433226 59832
rect 434720 59780 434772 59832
rect 435874 59780 435926 59832
rect 443000 59780 443052 59832
rect 443994 59780 444046 59832
rect 452660 59780 452712 59832
rect 453934 59780 453986 59832
rect 463792 59780 463844 59832
rect 464774 59780 464826 59832
rect 476212 59780 476264 59832
rect 477414 59780 477466 59832
rect 3424 59372 3476 59424
rect 69020 59372 69072 59424
rect 72424 57876 72476 57928
rect 85488 57876 85540 57928
rect 87604 57876 87656 57928
rect 92480 57876 92532 57928
rect 100668 57876 100720 57928
rect 57244 57808 57296 57860
rect 78312 57808 78364 57860
rect 88984 57808 89036 57860
rect 91836 57808 91888 57860
rect 97264 57808 97316 57860
rect 97908 57808 97960 57860
rect 98184 57808 98236 57860
rect 99196 57808 99248 57860
rect 99932 57808 99984 57860
rect 100576 57808 100628 57860
rect 100852 57808 100904 57860
rect 102048 57808 102100 57860
rect 109868 57876 109920 57928
rect 213736 57876 213788 57928
rect 305644 57876 305696 57928
rect 355508 57876 355560 57928
rect 358084 57876 358136 57928
rect 363604 57876 363656 57928
rect 364248 57876 364300 57928
rect 379888 57876 379940 57928
rect 392676 57876 392728 57928
rect 402428 57876 402480 57928
rect 155040 57808 155092 57860
rect 221832 57808 221884 57860
rect 322204 57808 322256 57860
rect 353668 57808 353720 57860
rect 378784 57808 378836 57860
rect 381544 57808 381596 57860
rect 400680 57808 400732 57860
rect 431224 57808 431276 57860
rect 437664 57876 437716 57928
rect 466368 57876 466420 57928
rect 484584 57876 484636 57928
rect 436744 57808 436796 57860
rect 438584 57808 438636 57860
rect 439504 57808 439556 57860
rect 440424 57808 440476 57860
rect 441528 57808 441580 57860
rect 478328 57808 478380 57860
rect 54484 57740 54536 57792
rect 114376 57740 114428 57792
rect 225512 57740 225564 57792
rect 340052 57740 340104 57792
rect 356428 57740 356480 57792
rect 357256 57740 357308 57792
rect 358268 57740 358320 57792
rect 358728 57740 358780 57792
rect 359096 57740 359148 57792
rect 360108 57740 360160 57792
rect 360936 57740 360988 57792
rect 361488 57740 361540 57792
rect 361856 57740 361908 57792
rect 362868 57740 362920 57792
rect 363604 57740 363656 57792
rect 451280 57740 451332 57792
rect 468392 57740 468444 57792
rect 483756 57740 483808 57792
rect 50344 57672 50396 57724
rect 106280 57672 106332 57724
rect 107108 57672 107160 57724
rect 115204 57672 115256 57724
rect 120724 57672 120776 57724
rect 155868 57672 155920 57724
rect 290464 57672 290516 57724
rect 298744 57672 298796 57724
rect 53104 57604 53156 57656
rect 113456 57604 113508 57656
rect 116584 57604 116636 57656
rect 117964 57604 118016 57656
rect 123484 57604 123536 57656
rect 124312 57604 124364 57656
rect 126244 57604 126296 57656
rect 127072 57604 127124 57656
rect 129740 57604 129792 57656
rect 130660 57604 130712 57656
rect 144184 57604 144236 57656
rect 145104 57604 145156 57656
rect 153200 57604 153252 57656
rect 154120 57604 154172 57656
rect 166264 57604 166316 57656
rect 167644 57604 167696 57656
rect 185768 57604 185820 57656
rect 186964 57604 187016 57656
rect 191196 57604 191248 57656
rect 191748 57604 191800 57656
rect 192024 57604 192076 57656
rect 193036 57604 193088 57656
rect 193864 57604 193916 57656
rect 194508 57604 194560 57656
rect 194784 57604 194836 57656
rect 195796 57604 195848 57656
rect 196624 57604 196676 57656
rect 197268 57604 197320 57656
rect 197452 57604 197504 57656
rect 198648 57604 198700 57656
rect 199292 57604 199344 57656
rect 200028 57604 200080 57656
rect 200212 57604 200264 57656
rect 201408 57604 201460 57656
rect 202052 57604 202104 57656
rect 202788 57604 202840 57656
rect 202880 57604 202932 57656
rect 204168 57604 204220 57656
rect 204720 57604 204772 57656
rect 205548 57604 205600 57656
rect 205640 57604 205692 57656
rect 206836 57604 206888 57656
rect 207388 57604 207440 57656
rect 208308 57604 208360 57656
rect 209228 57604 209280 57656
rect 209688 57604 209740 57656
rect 212816 57604 212868 57656
rect 213828 57604 213880 57656
rect 214656 57604 214708 57656
rect 215208 57604 215260 57656
rect 215576 57604 215628 57656
rect 216496 57604 216548 57656
rect 217324 57604 217376 57656
rect 217968 57604 218020 57656
rect 220084 57604 220136 57656
rect 220728 57604 220780 57656
rect 222752 57604 222804 57656
rect 223488 57604 223540 57656
rect 223672 57604 223724 57656
rect 224776 57604 224828 57656
rect 226432 57604 226484 57656
rect 227536 57604 227588 57656
rect 228180 57604 228232 57656
rect 229008 57604 229060 57656
rect 229100 57604 229152 57656
rect 230296 57604 230348 57656
rect 230940 57604 230992 57656
rect 231676 57604 231728 57656
rect 232688 57604 232740 57656
rect 233148 57604 233200 57656
rect 236368 57604 236420 57656
rect 238024 57604 238076 57656
rect 11704 57536 11756 57588
rect 71044 57536 71096 57588
rect 73804 57536 73856 57588
rect 79324 57536 79376 57588
rect 115940 57536 115992 57588
rect 124864 57536 124916 57588
rect 127900 57536 127952 57588
rect 129004 57536 129056 57588
rect 131580 57536 131632 57588
rect 148968 57536 149020 57588
rect 288440 57536 288492 57588
rect 289084 57536 289136 57588
rect 293960 57536 294012 57588
rect 299480 57536 299532 57588
rect 300400 57536 300452 57588
rect 306472 57672 306524 57724
rect 307668 57672 307720 57724
rect 331864 57672 331916 57724
rect 333796 57672 333848 57724
rect 343824 57672 343876 57724
rect 344928 57672 344980 57724
rect 345572 57672 345624 57724
rect 346308 57672 346360 57724
rect 346492 57672 346544 57724
rect 347688 57672 347740 57724
rect 348332 57672 348384 57724
rect 349068 57672 349120 57724
rect 349252 57672 349304 57724
rect 350356 57672 350408 57724
rect 351000 57672 351052 57724
rect 351828 57672 351880 57724
rect 351920 57672 351972 57724
rect 353208 57672 353260 57724
rect 353944 57672 353996 57724
rect 445760 57672 445812 57724
rect 458088 57672 458140 57724
rect 482836 57672 482888 57724
rect 364524 57604 364576 57656
rect 365536 57604 365588 57656
rect 366364 57604 366416 57656
rect 367008 57604 367060 57656
rect 367284 57604 367336 57656
rect 368388 57604 368440 57656
rect 369032 57604 369084 57656
rect 369768 57604 369820 57656
rect 369952 57604 370004 57656
rect 371148 57604 371200 57656
rect 371792 57604 371844 57656
rect 372528 57604 372580 57656
rect 372712 57604 372764 57656
rect 373908 57604 373960 57656
rect 374460 57604 374512 57656
rect 375288 57604 375340 57656
rect 375380 57604 375432 57656
rect 376576 57604 376628 57656
rect 377220 57604 377272 57656
rect 377956 57604 378008 57656
rect 378968 57604 379020 57656
rect 379428 57604 379480 57656
rect 381728 57604 381780 57656
rect 382188 57604 382240 57656
rect 382648 57604 382700 57656
rect 383476 57604 383528 57656
rect 418804 57604 418856 57656
rect 425060 57604 425112 57656
rect 425888 57604 425940 57656
rect 430488 57604 430540 57656
rect 317420 57536 317472 57588
rect 322940 57536 322992 57588
rect 323860 57536 323912 57588
rect 325700 57536 325752 57588
rect 326620 57536 326672 57588
rect 329932 57536 329984 57588
rect 331128 57536 331180 57588
rect 335360 57536 335412 57588
rect 336556 57536 336608 57588
rect 337476 57536 337528 57588
rect 338028 57536 338080 57588
rect 338396 57536 338448 57588
rect 339316 57536 339368 57588
rect 340144 57536 340196 57588
rect 340788 57536 340840 57588
rect 341064 57536 341116 57588
rect 342076 57536 342128 57588
rect 342904 57536 342956 57588
rect 343548 57536 343600 57588
rect 444840 57536 444892 57588
rect 448520 57536 448572 57588
rect 449348 57536 449400 57588
rect 471980 57604 472032 57656
rect 472900 57604 472952 57656
rect 480168 57604 480220 57656
rect 488264 57604 488316 57656
rect 491852 57604 491904 57656
rect 492864 57604 492916 57656
rect 494612 57604 494664 57656
rect 495348 57604 495400 57656
rect 495532 57604 495584 57656
rect 496728 57604 496780 57656
rect 497280 57604 497332 57656
rect 498108 57604 498160 57656
rect 498200 57604 498252 57656
rect 499396 57604 499448 57656
rect 500040 57604 500092 57656
rect 500776 57604 500828 57656
rect 501788 57604 501840 57656
rect 502248 57604 502300 57656
rect 505468 57604 505520 57656
rect 506388 57604 506440 57656
rect 507216 57604 507268 57656
rect 507768 57604 507820 57656
rect 508136 57604 508188 57656
rect 509056 57604 509108 57656
rect 509884 57604 509936 57656
rect 510528 57604 510580 57656
rect 510804 57604 510856 57656
rect 511816 57604 511868 57656
rect 513564 57604 513616 57656
rect 514576 57604 514628 57656
rect 515312 57604 515364 57656
rect 516048 57604 516100 57656
rect 516876 57604 516928 57656
rect 517428 57604 517480 57656
rect 475568 57536 475620 57588
rect 482928 57536 482980 57588
rect 489184 57536 489236 57588
rect 492772 57536 492824 57588
rect 493876 57536 493928 57588
rect 516232 57536 516284 57588
rect 517336 57536 517388 57588
rect 14464 57468 14516 57520
rect 75552 57468 75604 57520
rect 75828 57468 75880 57520
rect 148692 57468 148744 57520
rect 162124 57468 162176 57520
rect 171324 57468 171376 57520
rect 183008 57468 183060 57520
rect 184204 57468 184256 57520
rect 235448 57468 235500 57520
rect 384396 57468 384448 57520
rect 384948 57468 385000 57520
rect 385316 57468 385368 57520
rect 386328 57468 386380 57520
rect 387156 57468 387208 57520
rect 387708 57468 387760 57520
rect 387984 57468 388036 57520
rect 389088 57468 389140 57520
rect 389824 57468 389876 57520
rect 390468 57468 390520 57520
rect 390744 57468 390796 57520
rect 391848 57468 391900 57520
rect 392584 57468 392636 57520
rect 393228 57468 393280 57520
rect 393412 57468 393464 57520
rect 394608 57468 394660 57520
rect 395252 57468 395304 57520
rect 395988 57468 396040 57520
rect 396172 57468 396224 57520
rect 397276 57468 397328 57520
rect 398012 57468 398064 57520
rect 398748 57468 398800 57520
rect 400864 57468 400916 57520
rect 401600 57468 401652 57520
rect 401692 57468 401744 57520
rect 466552 57468 466604 57520
rect 467472 57468 467524 57520
rect 469128 57468 469180 57520
rect 485504 57468 485556 57520
rect 18604 57400 18656 57452
rect 134248 57400 134300 57452
rect 161388 57400 161440 57452
rect 176660 57400 176712 57452
rect 177304 57400 177356 57452
rect 179420 57400 179472 57452
rect 219164 57400 219216 57452
rect 222844 57400 222896 57452
rect 238116 57400 238168 57452
rect 238668 57400 238720 57452
rect 240876 57400 240928 57452
rect 241428 57400 241480 57452
rect 241704 57400 241756 57452
rect 242808 57400 242860 57452
rect 243544 57400 243596 57452
rect 244188 57400 244240 57452
rect 244464 57400 244516 57452
rect 245476 57400 245528 57452
rect 246212 57400 246264 57452
rect 246948 57400 247000 57452
rect 29644 57332 29696 57384
rect 164976 57332 165028 57384
rect 188436 57332 188488 57384
rect 196624 57332 196676 57384
rect 233608 57332 233660 57384
rect 239956 57332 240008 57384
rect 407764 57400 407816 57452
rect 410524 57400 410576 57452
rect 423220 57400 423272 57452
rect 423588 57400 423640 57452
rect 473820 57400 473872 57452
rect 476028 57400 476080 57452
rect 487344 57400 487396 57452
rect 512644 57400 512696 57452
rect 513288 57400 513340 57452
rect 247132 57332 247184 57384
rect 248328 57332 248380 57384
rect 248972 57332 249024 57384
rect 249708 57332 249760 57384
rect 249892 57332 249944 57384
rect 250996 57332 251048 57384
rect 251640 57332 251692 57384
rect 252468 57332 252520 57384
rect 252560 57332 252612 57384
rect 253756 57332 253808 57384
rect 254400 57332 254452 57384
rect 255228 57332 255280 57384
rect 255320 57332 255372 57384
rect 256608 57332 256660 57384
rect 257988 57332 258040 57384
rect 448428 57332 448480 57384
rect 455328 57332 455380 57384
rect 481916 57332 481968 57384
rect 22744 57264 22796 57316
rect 163136 57264 163188 57316
rect 165528 57264 165580 57316
rect 177580 57264 177632 57316
rect 190276 57264 190328 57316
rect 202144 57264 202196 57316
rect 208216 57264 208268 57316
rect 258724 57264 258776 57316
rect 258908 57264 258960 57316
rect 259368 57264 259420 57316
rect 261576 57264 261628 57316
rect 7564 57196 7616 57248
rect 166724 57196 166776 57248
rect 183928 57196 183980 57248
rect 188436 57196 188488 57248
rect 189356 57196 189408 57248
rect 204904 57196 204956 57248
rect 210148 57196 210200 57248
rect 264244 57196 264296 57248
rect 489184 57264 489236 57316
rect 265256 57196 265308 57248
rect 507124 57196 507176 57248
rect 68284 57128 68336 57180
rect 84568 57128 84620 57180
rect 211988 57128 212040 57180
rect 69664 57060 69716 57112
rect 83648 57060 83700 57112
rect 257068 57060 257120 57112
rect 257988 57060 258040 57112
rect 262864 57060 262916 57112
rect 287704 57128 287756 57180
rect 293224 57128 293276 57180
rect 342904 57128 342956 57180
rect 371884 57128 371936 57180
rect 389824 57128 389876 57180
rect 450544 57128 450596 57180
rect 462228 57128 462280 57180
rect 473268 57128 473320 57180
rect 486424 57128 486476 57180
rect 504548 57128 504600 57180
rect 505008 57128 505060 57180
rect 315764 57060 315816 57112
rect 480076 57060 480128 57112
rect 71780 56992 71832 57044
rect 81900 56992 81952 57044
rect 239036 56992 239088 57044
rect 246304 56992 246356 57044
rect 264336 56992 264388 57044
rect 264888 56992 264940 57044
rect 267004 56992 267056 57044
rect 267648 56992 267700 57044
rect 267924 56992 267976 57044
rect 269028 56992 269080 57044
rect 269764 56992 269816 57044
rect 270408 56992 270460 57044
rect 270684 56992 270736 57044
rect 271696 56992 271748 57044
rect 272432 56992 272484 57044
rect 273168 56992 273220 57044
rect 65616 56924 65668 56976
rect 278136 56924 278188 56976
rect 320180 56992 320232 57044
rect 502708 56992 502760 57044
rect 503536 56992 503588 57044
rect 284944 56856 284996 56908
rect 316684 56856 316736 56908
rect 319352 56856 319404 56908
rect 86224 56788 86276 56840
rect 89996 56788 90048 56840
rect 186688 56720 186740 56772
rect 191104 56720 191156 56772
rect 221004 56720 221056 56772
rect 228364 56720 228416 56772
rect 237196 56652 237248 56704
rect 240784 56652 240836 56704
rect 373632 56652 373684 56704
rect 374644 56652 374696 56704
rect 102692 56584 102744 56636
rect 105544 56584 105596 56636
rect 170404 56584 170456 56636
rect 172152 56584 172204 56636
rect 179328 56584 179380 56636
rect 181260 56584 181312 56636
rect 218244 56584 218296 56636
rect 220084 56584 220136 56636
rect 273352 56584 273404 56636
rect 274456 56584 274508 56636
rect 275192 56584 275244 56636
rect 275928 56584 275980 56636
rect 276020 56584 276072 56636
rect 277308 56584 277360 56636
rect 277860 56584 277912 56636
rect 278688 56584 278740 56636
rect 278780 56584 278832 56636
rect 280068 56584 280120 56636
rect 280528 56584 280580 56636
rect 281356 56584 281408 56636
rect 282368 56584 282420 56636
rect 282828 56584 282880 56636
rect 295984 56584 296036 56636
rect 296812 56584 296864 56636
rect 421564 56584 421616 56636
rect 422300 56584 422352 56636
rect 487068 56584 487120 56636
rect 490012 56584 490064 56636
rect 62028 56380 62080 56432
rect 87328 56380 87380 56432
rect 41328 56312 41380 56364
rect 71780 56312 71832 56364
rect 37188 56244 37240 56296
rect 80980 56244 81032 56296
rect 345664 56244 345716 56296
rect 452108 56244 452160 56296
rect 34428 56176 34480 56228
rect 79968 56176 80020 56228
rect 188344 56176 188396 56228
rect 297732 56176 297784 56228
rect 380808 56176 380860 56228
rect 501604 56176 501656 56228
rect 22008 56108 22060 56160
rect 77208 56108 77260 56160
rect 282184 56108 282236 56160
rect 434076 56108 434128 56160
rect 43444 56040 43496 56092
rect 109040 56040 109092 56092
rect 260104 56040 260156 56092
rect 427728 56040 427780 56092
rect 25504 55972 25556 56024
rect 103520 55972 103572 56024
rect 249064 55972 249116 56024
rect 426808 55972 426860 56024
rect 65524 55904 65576 55956
rect 146024 55904 146076 55956
rect 262496 55904 262548 55956
rect 483664 55904 483716 55956
rect 58624 55836 58676 55888
rect 142344 55836 142396 55888
rect 259828 55836 259880 55888
rect 485044 55836 485096 55888
rect 47584 54680 47636 54732
rect 110512 54680 110564 54732
rect 39304 54612 39356 54664
rect 106372 54612 106424 54664
rect 35164 54544 35216 54596
rect 104900 54544 104952 54596
rect 318064 54544 318116 54596
rect 440516 54544 440568 54596
rect 15844 54476 15896 54528
rect 132592 54476 132644 54528
rect 251824 54476 251876 54528
rect 429292 54476 429344 54528
rect 519820 46860 519872 46912
rect 580172 46860 580224 46912
rect 267004 37884 267056 37936
rect 429200 37884 429252 37936
rect 142068 36524 142120 36576
rect 285772 36524 285824 36576
rect 286324 36524 286376 36576
rect 432052 36524 432104 36576
rect 233884 33736 233936 33788
rect 425152 33736 425204 33788
rect 519728 33056 519780 33108
rect 580172 33056 580224 33108
rect 160008 32376 160060 32428
rect 291292 32376 291344 32428
rect 360844 32376 360896 32428
rect 449900 32376 449952 32428
rect 153108 31016 153160 31068
rect 288532 31016 288584 31068
rect 320824 31016 320876 31068
rect 443092 31016 443144 31068
rect 61936 29588 61988 29640
rect 144184 29588 144236 29640
rect 209044 29588 209096 29640
rect 299572 29588 299624 29640
rect 374644 29588 374696 29640
rect 481640 29588 481692 29640
rect 144828 28228 144880 28280
rect 170404 28228 170456 28280
rect 289176 28228 289228 28280
rect 434812 28228 434864 28280
rect 173808 26868 173860 26920
rect 294052 26868 294104 26920
rect 300124 26868 300176 26920
rect 441620 26868 441672 26920
rect 51724 25508 51776 25560
rect 111800 25508 111852 25560
rect 113088 25508 113140 25560
rect 129832 25508 129884 25560
rect 222844 25508 222896 25560
rect 327172 25508 327224 25560
rect 376576 25508 376628 25560
rect 486424 25508 486476 25560
rect 81348 24080 81400 24132
rect 121460 24080 121512 24132
rect 241428 24080 241480 24132
rect 412732 24080 412784 24132
rect 376024 22788 376076 22840
rect 452752 22788 452804 22840
rect 238024 22720 238076 22772
rect 394700 22720 394752 22772
rect 224776 21428 224828 21480
rect 345020 21428 345072 21480
rect 238024 21360 238076 21412
rect 423680 21360 423732 21412
rect 519636 20612 519688 20664
rect 579988 20612 580040 20664
rect 228364 20000 228416 20052
rect 334072 20000 334124 20052
rect 374644 20000 374696 20052
rect 454040 20000 454092 20052
rect 59268 19932 59320 19984
rect 85580 19932 85632 19984
rect 224776 19932 224828 19984
rect 410524 19932 410576 19984
rect 220084 18640 220136 18692
rect 324412 18640 324464 18692
rect 68376 18572 68428 18624
rect 143540 18572 143592 18624
rect 220636 18572 220688 18624
rect 421564 18572 421616 18624
rect 358084 17484 358136 17536
rect 409972 17484 410024 17536
rect 216496 17416 216548 17468
rect 313372 17416 313424 17468
rect 358176 17416 358228 17468
rect 448612 17416 448664 17468
rect 294604 17348 294656 17400
rect 438860 17348 438912 17400
rect 269764 17280 269816 17332
rect 430580 17280 430632 17332
rect 32404 17212 32456 17264
rect 78680 17212 78732 17264
rect 143448 17212 143500 17264
rect 392584 17212 392636 17264
rect 211068 16260 211120 16312
rect 295616 16260 295668 16312
rect 377956 16192 378008 16244
rect 468484 16192 468536 16244
rect 180064 16124 180116 16176
rect 295432 16124 295484 16176
rect 323584 16124 323636 16176
rect 447140 16124 447192 16176
rect 291844 16056 291896 16108
rect 436100 16056 436152 16108
rect 240876 15988 240928 16040
rect 425060 15988 425112 16040
rect 220084 15920 220136 15972
rect 420920 15920 420972 15972
rect 52368 15852 52420 15904
rect 68284 15852 68336 15904
rect 139308 15852 139360 15904
rect 400864 15852 400916 15904
rect 259276 14900 259328 14952
rect 316040 14900 316092 14952
rect 169576 14832 169628 14884
rect 289084 14832 289136 14884
rect 377404 14832 377456 14884
rect 452660 14832 452712 14884
rect 144736 14764 144788 14816
rect 287060 14764 287112 14816
rect 287796 14764 287848 14816
rect 434720 14764 434772 14816
rect 137652 14696 137704 14748
rect 285680 14696 285732 14748
rect 292488 14696 292540 14748
rect 439504 14696 439556 14748
rect 240784 14628 240836 14680
rect 398840 14628 398892 14680
rect 246304 14560 246356 14612
rect 406016 14560 406068 14612
rect 246396 14492 246448 14544
rect 427820 14492 427872 14544
rect 54944 14424 54996 14476
rect 65616 14424 65668 14476
rect 259368 14424 259420 14476
rect 483664 14424 483716 14476
rect 268844 13676 268896 13728
rect 316684 13676 316736 13728
rect 216588 13608 216640 13660
rect 316040 13608 316092 13660
rect 220728 13540 220780 13592
rect 331588 13540 331640 13592
rect 379428 13540 379480 13592
rect 471244 13540 471296 13592
rect 224868 13472 224920 13524
rect 349252 13472 349304 13524
rect 353944 13472 353996 13524
rect 448520 13472 448572 13524
rect 180708 13404 180760 13456
rect 295984 13404 296036 13456
rect 316776 13404 316828 13456
rect 443000 13404 443052 13456
rect 227536 13336 227588 13388
rect 356336 13336 356388 13388
rect 378048 13336 378100 13388
rect 497464 13336 497516 13388
rect 281264 13268 281316 13320
rect 431224 13268 431276 13320
rect 234528 13200 234580 13252
rect 387800 13200 387852 13252
rect 264336 13132 264388 13184
rect 431960 13132 432012 13184
rect 17868 13064 17920 13116
rect 75920 13064 75972 13116
rect 76564 13064 76616 13116
rect 147772 13064 147824 13116
rect 202144 13064 202196 13116
rect 214472 13064 214524 13116
rect 264888 13064 264940 13116
rect 504364 13064 504416 13116
rect 209688 12384 209740 12436
rect 288992 12384 289044 12436
rect 213828 12316 213880 12368
rect 303160 12316 303212 12368
rect 378784 12316 378836 12368
rect 403624 12316 403676 12368
rect 215208 12248 215260 12300
rect 309784 12248 309836 12300
rect 354588 12248 354640 12300
rect 407120 12248 407172 12300
rect 223488 12180 223540 12232
rect 340880 12180 340932 12232
rect 375288 12180 375340 12232
rect 484768 12180 484820 12232
rect 217968 12112 218020 12164
rect 320456 12112 320508 12164
rect 322296 12112 322348 12164
rect 445852 12112 445904 12164
rect 227628 12044 227680 12096
rect 359464 12044 359516 12096
rect 376668 12044 376720 12096
rect 490564 12044 490616 12096
rect 285588 11976 285640 12028
rect 436744 11976 436796 12028
rect 238668 11908 238720 11960
rect 402520 11908 402572 11960
rect 260656 11840 260708 11892
rect 489276 11840 489328 11892
rect 57336 11772 57388 11824
rect 142160 11772 142212 11824
rect 263416 11772 263468 11824
rect 501328 11772 501380 11824
rect 136456 11704 136508 11756
rect 381544 11704 381596 11756
rect 192944 10956 192996 11008
rect 414020 10956 414072 11008
rect 188988 10888 189040 10940
rect 414112 10888 414164 10940
rect 186228 10820 186280 10872
rect 412640 10820 412692 10872
rect 182088 10752 182140 10804
rect 411260 10752 411312 10804
rect 177856 10684 177908 10736
rect 411352 10684 411404 10736
rect 175188 10616 175240 10668
rect 409880 10616 409932 10668
rect 170772 10548 170824 10600
rect 408592 10548 408644 10600
rect 168288 10480 168340 10532
rect 408500 10480 408552 10532
rect 164148 10412 164200 10464
rect 407212 10412 407264 10464
rect 131764 10344 131816 10396
rect 399024 10344 399076 10396
rect 66168 10276 66220 10328
rect 86960 10276 87012 10328
rect 128176 10276 128228 10328
rect 398932 10276 398984 10328
rect 418804 10276 418856 10328
rect 506480 10276 506532 10328
rect 195612 10208 195664 10260
rect 415400 10208 415452 10260
rect 199936 10140 199988 10192
rect 416872 10140 416924 10192
rect 202696 10072 202748 10124
rect 416780 10072 416832 10124
rect 206744 10004 206796 10056
rect 418160 10004 418212 10056
rect 211068 9936 211120 9988
rect 419632 9936 419684 9988
rect 213828 9868 213880 9920
rect 419540 9868 419592 9920
rect 277124 9800 277176 9852
rect 320272 9800 320324 9852
rect 279516 9732 279568 9784
rect 321560 9732 321612 9784
rect 222752 9596 222804 9648
rect 306472 9596 306524 9648
rect 364248 9596 364300 9648
rect 442632 9596 442684 9648
rect 219256 9528 219308 9580
rect 306380 9528 306432 9580
rect 365536 9528 365588 9580
rect 446220 9528 446272 9580
rect 215668 9460 215720 9512
rect 305000 9460 305052 9512
rect 365628 9460 365680 9512
rect 449808 9460 449860 9512
rect 212172 9392 212224 9444
rect 303620 9392 303672 9444
rect 367008 9392 367060 9444
rect 453304 9392 453356 9444
rect 208584 9324 208636 9376
rect 303712 9324 303764 9376
rect 368388 9324 368440 9376
rect 456892 9324 456944 9376
rect 205088 9256 205140 9308
rect 302424 9256 302476 9308
rect 368296 9256 368348 9308
rect 460388 9256 460440 9308
rect 201500 9188 201552 9240
rect 302332 9188 302384 9240
rect 369768 9188 369820 9240
rect 463976 9188 464028 9240
rect 197912 9120 197964 9172
rect 300860 9120 300912 9172
rect 371148 9120 371200 9172
rect 467472 9120 467524 9172
rect 194416 9052 194468 9104
rect 299480 9052 299532 9104
rect 325608 9052 325660 9104
rect 331864 9052 331916 9104
rect 371056 9052 371108 9104
rect 471060 9052 471112 9104
rect 47860 8916 47912 8968
rect 69664 8984 69716 9036
rect 134156 8984 134208 9036
rect 284300 8984 284352 9036
rect 322204 8984 322256 9036
rect 338672 8984 338724 9036
rect 340144 8984 340196 9036
rect 352840 8984 352892 9036
rect 372528 8984 372580 9036
rect 474556 8984 474608 9036
rect 69112 8916 69164 8968
rect 88340 8916 88392 8968
rect 105728 8916 105780 8968
rect 124864 8916 124916 8968
rect 130568 8916 130620 8968
rect 283012 8916 283064 8968
rect 312636 8916 312688 8968
rect 353852 8916 353904 8968
rect 373908 8916 373960 8968
rect 478144 8916 478196 8968
rect 226340 8848 226392 8900
rect 307760 8848 307812 8900
rect 362776 8848 362828 8900
rect 439136 8848 439188 8900
rect 229836 8780 229888 8832
rect 309232 8780 309284 8832
rect 362868 8780 362920 8832
rect 435548 8780 435600 8832
rect 233424 8712 233476 8764
rect 309324 8712 309376 8764
rect 361488 8712 361540 8764
rect 432052 8712 432104 8764
rect 237012 8644 237064 8696
rect 310520 8644 310572 8696
rect 360016 8644 360068 8696
rect 428464 8644 428516 8696
rect 240508 8576 240560 8628
rect 311900 8576 311952 8628
rect 360108 8576 360160 8628
rect 424968 8576 425020 8628
rect 244096 8508 244148 8560
rect 311992 8508 312044 8560
rect 358728 8508 358780 8560
rect 421380 8508 421432 8560
rect 247592 8440 247644 8492
rect 313280 8440 313332 8492
rect 357348 8440 357400 8492
rect 417884 8440 417936 8492
rect 251180 8372 251232 8424
rect 314752 8372 314804 8424
rect 357256 8372 357308 8424
rect 414296 8372 414348 8424
rect 305644 8304 305696 8356
rect 306748 8304 306800 8356
rect 52552 8236 52604 8288
rect 54484 8236 54536 8288
rect 248236 8236 248288 8288
rect 441252 8236 441304 8288
rect 249708 8168 249760 8220
rect 445024 8168 445076 8220
rect 250996 8100 251048 8152
rect 448612 8100 448664 8152
rect 450544 8100 450596 8152
rect 480536 8100 480588 8152
rect 251088 8032 251140 8084
rect 452108 8032 452160 8084
rect 252468 7964 252520 8016
rect 455696 7964 455748 8016
rect 253756 7896 253808 7948
rect 459192 7896 459244 7948
rect 253848 7828 253900 7880
rect 462780 7828 462832 7880
rect 255228 7760 255280 7812
rect 466276 7760 466328 7812
rect 256608 7692 256660 7744
rect 469864 7692 469916 7744
rect 70308 7624 70360 7676
rect 118700 7624 118752 7676
rect 256516 7624 256568 7676
rect 473452 7624 473504 7676
rect 42984 7556 43036 7608
rect 110420 7556 110472 7608
rect 119896 7556 119948 7608
rect 129004 7556 129056 7608
rect 257988 7556 258040 7608
rect 476948 7556 477000 7608
rect 248328 7488 248380 7540
rect 437940 7488 437992 7540
rect 246948 7420 247000 7472
rect 434444 7420 434496 7472
rect 245568 7352 245620 7404
rect 430856 7352 430908 7404
rect 245476 7284 245528 7336
rect 427268 7284 427320 7336
rect 244188 7216 244240 7268
rect 423772 7216 423824 7268
rect 242716 7148 242768 7200
rect 420184 7148 420236 7200
rect 242808 7080 242860 7132
rect 416688 7080 416740 7132
rect 126980 7012 127032 7064
rect 282920 7012 282972 7064
rect 283104 7012 283156 7064
rect 323032 7012 323084 7064
rect 353116 7012 353168 7064
rect 400128 7012 400180 7064
rect 261760 6808 261812 6860
rect 298744 6808 298796 6860
rect 304356 6808 304408 6860
rect 328460 6808 328512 6860
rect 347596 6808 347648 6860
rect 378876 6808 378928 6860
rect 389824 6808 389876 6860
rect 391848 6808 391900 6860
rect 519544 6808 519596 6860
rect 580172 6808 580224 6860
rect 265348 6740 265400 6792
rect 317512 6740 317564 6792
rect 318524 6740 318576 6792
rect 331220 6740 331272 6792
rect 349068 6740 349120 6792
rect 382372 6740 382424 6792
rect 390468 6740 390520 6792
rect 545488 6740 545540 6792
rect 187332 6672 187384 6724
rect 298100 6672 298152 6724
rect 300768 6672 300820 6724
rect 327080 6672 327132 6724
rect 350356 6672 350408 6724
rect 385960 6672 386012 6724
rect 391756 6672 391808 6724
rect 549076 6672 549128 6724
rect 102232 6604 102284 6656
rect 126244 6604 126296 6656
rect 166080 6604 166132 6656
rect 287704 6604 287756 6656
rect 290188 6604 290240 6656
rect 324320 6604 324372 6656
rect 350448 6604 350500 6656
rect 389456 6604 389508 6656
rect 391664 6604 391716 6656
rect 552664 6604 552716 6656
rect 98644 6536 98696 6588
rect 125600 6536 125652 6588
rect 162492 6536 162544 6588
rect 291200 6536 291252 6588
rect 293684 6536 293736 6588
rect 325792 6536 325844 6588
rect 340788 6536 340840 6588
rect 350356 6536 350408 6588
rect 351828 6536 351880 6588
rect 393044 6536 393096 6588
rect 393228 6536 393280 6588
rect 556160 6536 556212 6588
rect 95056 6468 95108 6520
rect 124312 6468 124364 6520
rect 229008 6468 229060 6520
rect 363512 6468 363564 6520
rect 394608 6468 394660 6520
rect 559748 6468 559800 6520
rect 87972 6400 88024 6452
rect 122840 6400 122892 6452
rect 230296 6400 230348 6452
rect 367008 6400 367060 6452
rect 394516 6400 394568 6452
rect 563244 6400 563296 6452
rect 63224 6332 63276 6384
rect 116032 6332 116084 6384
rect 230388 6332 230440 6384
rect 370596 6332 370648 6384
rect 371884 6332 371936 6384
rect 384764 6332 384816 6384
rect 395988 6332 396040 6384
rect 566832 6332 566884 6384
rect 2872 6264 2924 6316
rect 71044 6264 71096 6316
rect 71228 6264 71280 6316
rect 146300 6264 146352 6316
rect 231676 6264 231728 6316
rect 374092 6264 374144 6316
rect 396540 6264 396592 6316
rect 397276 6264 397328 6316
rect 570328 6264 570380 6316
rect 27712 6196 27764 6248
rect 107660 6196 107712 6248
rect 116400 6196 116452 6248
rect 129740 6196 129792 6248
rect 196624 6196 196676 6248
rect 207388 6196 207440 6248
rect 231768 6196 231820 6248
rect 377680 6196 377732 6248
rect 388996 6196 389048 6248
rect 397368 6196 397420 6248
rect 573916 6196 573968 6248
rect 23020 6128 23072 6180
rect 106280 6128 106332 6180
rect 125876 6128 125928 6180
rect 166264 6128 166316 6180
rect 186964 6128 187016 6180
rect 196808 6128 196860 6180
rect 233148 6128 233200 6180
rect 381176 6128 381228 6180
rect 387708 6128 387760 6180
rect 258724 6060 258776 6112
rect 285404 6060 285456 6112
rect 286600 6060 286652 6112
rect 322940 6060 322992 6112
rect 342076 6060 342128 6112
rect 347688 6060 347740 6112
rect 375288 6060 375340 6112
rect 389088 6060 389140 6112
rect 264244 5992 264296 6044
rect 292580 5992 292632 6044
rect 297272 5992 297324 6044
rect 325700 5992 325752 6044
rect 346308 5992 346360 6044
rect 371700 5992 371752 6044
rect 384948 5992 385000 6044
rect 398748 6128 398800 6180
rect 577412 6128 577464 6180
rect 538404 6060 538456 6112
rect 534908 5992 534960 6044
rect 284944 5924 284996 5976
rect 299664 5924 299716 5976
rect 307944 5924 307996 5976
rect 328552 5924 328604 5976
rect 344836 5924 344888 5976
rect 368204 5924 368256 5976
rect 386236 5924 386288 5976
rect 531320 5924 531372 5976
rect 311440 5856 311492 5908
rect 329840 5856 329892 5908
rect 344928 5856 344980 5908
rect 364616 5856 364668 5908
rect 386328 5856 386380 5908
rect 527824 5856 527876 5908
rect 315028 5788 315080 5840
rect 329932 5788 329984 5840
rect 343548 5788 343600 5840
rect 361120 5788 361172 5840
rect 524236 5788 524288 5840
rect 322112 5720 322164 5772
rect 332692 5720 332744 5772
rect 342168 5720 342220 5772
rect 357532 5720 357584 5772
rect 383568 5720 383620 5772
rect 520740 5720 520792 5772
rect 339408 5652 339460 5704
rect 346952 5652 347004 5704
rect 354036 5652 354088 5704
rect 383476 5652 383528 5704
rect 517152 5652 517204 5704
rect 332692 5584 332744 5636
rect 335452 5584 335504 5636
rect 339316 5584 339368 5636
rect 343364 5584 343416 5636
rect 382188 5584 382240 5636
rect 513564 5584 513616 5636
rect 204904 5516 204956 5568
rect 210976 5516 211028 5568
rect 329196 5516 329248 5568
rect 333980 5516 334032 5568
rect 338028 5516 338080 5568
rect 339868 5516 339920 5568
rect 353208 5516 353260 5568
rect 541992 5516 542044 5568
rect 100576 5448 100628 5500
rect 111616 5448 111668 5500
rect 198556 5448 198608 5500
rect 246304 5448 246356 5500
rect 274456 5448 274508 5500
rect 540796 5448 540848 5500
rect 83280 5380 83332 5432
rect 87604 5380 87656 5432
rect 102048 5380 102100 5432
rect 115112 5380 115164 5432
rect 200028 5380 200080 5432
rect 249984 5380 250036 5432
rect 274548 5380 274600 5432
rect 544384 5380 544436 5432
rect 76196 5312 76248 5364
rect 89812 5312 89864 5364
rect 105544 5312 105596 5364
rect 122288 5312 122340 5364
rect 201408 5312 201460 5364
rect 253480 5312 253532 5364
rect 254676 5312 254728 5364
rect 262864 5312 262916 5364
rect 275928 5312 275980 5364
rect 547880 5312 547932 5364
rect 72608 5244 72660 5296
rect 86224 5244 86276 5296
rect 101956 5244 102008 5296
rect 118792 5244 118844 5296
rect 201316 5244 201368 5296
rect 257068 5244 257120 5296
rect 277308 5244 277360 5296
rect 551468 5244 551520 5296
rect 59636 5176 59688 5228
rect 79324 5176 79376 5228
rect 79692 5176 79744 5228
rect 88984 5176 89036 5228
rect 91560 5176 91612 5228
rect 123484 5176 123536 5228
rect 202788 5176 202840 5228
rect 260656 5176 260708 5228
rect 277216 5176 277268 5228
rect 554964 5176 555016 5228
rect 44272 5108 44324 5160
rect 82820 5108 82872 5160
rect 84476 5108 84528 5160
rect 121644 5108 121696 5160
rect 204168 5108 204220 5160
rect 264152 5108 264204 5160
rect 279976 5108 280028 5160
rect 558552 5108 558604 5160
rect 26516 5040 26568 5092
rect 57244 5040 57296 5092
rect 66720 5040 66772 5092
rect 116584 5040 116636 5092
rect 140044 5040 140096 5092
rect 162124 5040 162176 5092
rect 204076 5040 204128 5092
rect 267740 5040 267792 5092
rect 280068 5040 280120 5092
rect 562048 5040 562100 5092
rect 34796 4972 34848 5024
rect 50344 4972 50396 5024
rect 56048 4972 56100 5024
rect 114652 4972 114704 5024
rect 147128 4972 147180 5024
rect 172520 4972 172572 5024
rect 205548 4972 205600 5024
rect 271236 4972 271288 5024
rect 271696 4972 271748 5024
rect 565636 4972 565688 5024
rect 7656 4904 7708 4956
rect 74632 4904 74684 4956
rect 77392 4904 77444 4956
rect 115204 4904 115256 4956
rect 136548 4904 136600 4956
rect 169760 4904 169812 4956
rect 184848 4904 184900 4956
rect 193220 4904 193272 4956
rect 206836 4904 206888 4956
rect 274824 4904 274876 4956
rect 281356 4904 281408 4956
rect 569132 4904 569184 4956
rect 572 4836 624 4888
rect 71872 4836 71924 4888
rect 73804 4836 73856 4888
rect 118884 4836 118936 4888
rect 123484 4836 123536 4888
rect 132500 4836 132552 4888
rect 132960 4836 133012 4888
rect 168380 4836 168432 4888
rect 191104 4836 191156 4888
rect 200304 4836 200356 4888
rect 206928 4836 206980 4888
rect 272616 4836 272668 4888
rect 278044 4836 278096 4888
rect 281448 4836 281500 4888
rect 572720 4836 572772 4888
rect 8760 4768 8812 4820
rect 103704 4768 103756 4820
rect 109316 4768 109368 4820
rect 128360 4768 128412 4820
rect 129372 4768 129424 4820
rect 168472 4768 168524 4820
rect 187608 4768 187660 4820
rect 203892 4768 203944 4820
rect 208308 4768 208360 4820
rect 281908 4768 281960 4820
rect 282828 4768 282880 4820
rect 576308 4768 576360 4820
rect 99288 4700 99340 4752
rect 108120 4700 108172 4752
rect 198648 4700 198700 4752
rect 242900 4700 242952 4752
rect 278320 4700 278372 4752
rect 197268 4632 197320 4684
rect 239312 4632 239364 4684
rect 273168 4632 273220 4684
rect 537208 4700 537260 4752
rect 99196 4564 99248 4616
rect 104532 4564 104584 4616
rect 195888 4564 195940 4616
rect 235816 4564 235868 4616
rect 271788 4564 271840 4616
rect 533712 4632 533764 4684
rect 530124 4564 530176 4616
rect 90364 4496 90416 4548
rect 93860 4496 93912 4548
rect 195796 4496 195848 4548
rect 232228 4496 232280 4548
rect 270408 4496 270460 4548
rect 526628 4496 526680 4548
rect 194508 4428 194560 4480
rect 228732 4428 228784 4480
rect 268936 4428 268988 4480
rect 523040 4428 523092 4480
rect 193128 4360 193180 4412
rect 225144 4360 225196 4412
rect 269028 4360 269080 4412
rect 519544 4360 519596 4412
rect 193036 4292 193088 4344
rect 221556 4292 221608 4344
rect 267648 4292 267700 4344
rect 515956 4292 516008 4344
rect 191748 4224 191800 4276
rect 218060 4224 218112 4276
rect 266268 4224 266320 4276
rect 512460 4224 512512 4276
rect 48964 4156 49016 4208
rect 53104 4156 53156 4208
rect 86868 4156 86920 4208
rect 92572 4156 92624 4208
rect 97908 4156 97960 4208
rect 101036 4156 101088 4208
rect 188436 4156 188488 4208
rect 189724 4156 189776 4208
rect 278688 4156 278740 4208
rect 407764 4156 407816 4208
rect 409604 4156 409656 4208
rect 53748 4088 53800 4140
rect 57336 4088 57388 4140
rect 64328 4088 64380 4140
rect 65432 4088 65484 4140
rect 71504 4088 71556 4140
rect 76564 4088 76616 4140
rect 89168 4088 89220 4140
rect 45468 4020 45520 4072
rect 51724 4020 51776 4072
rect 85672 4020 85724 4072
rect 150440 4020 150492 4072
rect 234620 4088 234672 4140
rect 240876 4088 240928 4140
rect 344560 4088 344612 4140
rect 377404 4088 377456 4140
rect 383568 4088 383620 4140
rect 463884 4088 463936 4140
rect 489276 4088 489328 4140
rect 491116 4088 491168 4140
rect 506296 4088 506348 4140
rect 550272 4088 550324 4140
rect 255872 4020 255924 4072
rect 269764 4020 269816 4072
rect 273628 4020 273680 4072
rect 287796 4020 287848 4072
rect 340972 4020 341024 4072
rect 376024 4020 376076 4072
rect 379980 4020 380032 4072
rect 462320 4020 462372 4072
rect 507768 4020 507820 4072
rect 553768 4020 553820 4072
rect 14740 3952 14792 4004
rect 18604 3952 18656 4004
rect 50160 3952 50212 4004
rect 58624 3952 58676 4004
rect 82084 3952 82136 4004
rect 150532 3952 150584 4004
rect 151820 3952 151872 4004
rect 160376 3952 160428 4004
rect 168380 3952 168432 4004
rect 178040 3952 178092 4004
rect 216864 3952 216916 4004
rect 220084 3952 220136 4004
rect 266544 3952 266596 4004
rect 282184 3952 282236 4004
rect 305552 3952 305604 4004
rect 316776 3952 316828 4004
rect 333888 3952 333940 4004
rect 363604 3952 363656 4004
rect 376484 3952 376536 4004
rect 461032 3952 461084 4004
rect 509056 3952 509108 4004
rect 557356 3952 557408 4004
rect 38384 3884 38436 3936
rect 47584 3884 47636 3936
rect 57244 3884 57296 3936
rect 68376 3884 68428 3936
rect 78588 3884 78640 3936
rect 149060 3884 149112 3936
rect 157800 3884 157852 3936
rect 175280 3884 175332 3936
rect 252376 3884 252428 3936
rect 267004 3884 267056 3936
rect 277216 3884 277268 3936
rect 291844 3884 291896 3936
rect 301964 3884 302016 3936
rect 320824 3884 320876 3936
rect 330392 3884 330444 3936
rect 360844 3884 360896 3936
rect 372896 3884 372948 3936
rect 460940 3884 460992 3936
rect 509148 3884 509200 3936
rect 560852 3884 560904 3936
rect 31300 3816 31352 3868
rect 43444 3816 43496 3868
rect 46664 3816 46716 3868
rect 140780 3816 140832 3868
rect 154212 3816 154264 3868
rect 173900 3816 173952 3868
rect 227536 3816 227588 3868
rect 238024 3816 238076 3868
rect 241704 3816 241756 3868
rect 260104 3816 260156 3868
rect 270040 3816 270092 3868
rect 289176 3816 289228 3868
rect 309048 3816 309100 3868
rect 342904 3816 342956 3868
rect 369400 3816 369452 3868
rect 18236 3748 18288 3800
rect 39304 3748 39356 3800
rect 43076 3748 43128 3800
rect 139400 3748 139452 3800
rect 150624 3748 150676 3800
rect 173992 3748 174044 3800
rect 190828 3748 190880 3800
rect 209044 3748 209096 3800
rect 238116 3748 238168 3800
rect 249064 3748 249116 3800
rect 259460 3748 259512 3800
rect 286324 3748 286376 3800
rect 294880 3748 294932 3800
rect 318064 3748 318116 3800
rect 323308 3748 323360 3800
rect 358176 3748 358228 3800
rect 365812 3748 365864 3800
rect 458364 3816 458416 3868
rect 472072 3816 472124 3868
rect 495348 3816 495400 3868
rect 504180 3816 504232 3868
rect 510528 3816 510580 3868
rect 564440 3816 564492 3868
rect 39580 3680 39632 3732
rect 136824 3680 136876 3732
rect 160100 3680 160152 3732
rect 405740 3680 405792 3732
rect 418988 3680 419040 3732
rect 454500 3680 454552 3732
rect 455328 3680 455380 3732
rect 459560 3680 459612 3732
rect 468484 3748 468536 3800
rect 495900 3748 495952 3800
rect 496636 3748 496688 3800
rect 511816 3748 511868 3800
rect 568028 3748 568080 3800
rect 471980 3680 472032 3732
rect 496728 3680 496780 3732
rect 507676 3680 507728 3732
rect 511908 3680 511960 3732
rect 571524 3680 571576 3732
rect 13544 3612 13596 3664
rect 35164 3612 35216 3664
rect 35992 3612 36044 3664
rect 138020 3612 138072 3664
rect 156604 3612 156656 3664
rect 405832 3612 405884 3664
rect 422576 3612 422628 3664
rect 423588 3612 423640 3664
rect 429660 3612 429712 3664
rect 430488 3612 430540 3664
rect 469312 3612 469364 3664
rect 486424 3612 486476 3664
rect 488816 3612 488868 3664
rect 489184 3612 489236 3664
rect 494704 3612 494756 3664
rect 498108 3612 498160 3664
rect 9956 3544 10008 3596
rect 15844 3544 15896 3596
rect 25320 3544 25372 3596
rect 29644 3544 29696 3596
rect 32496 3544 32548 3596
rect 136640 3544 136692 3596
rect 151820 3544 151872 3596
rect 153108 3544 153160 3596
rect 155408 3544 155460 3596
rect 155868 3544 155920 3596
rect 158904 3544 158956 3596
rect 160008 3544 160060 3596
rect 404360 3544 404412 3596
rect 411904 3544 411956 3596
rect 470600 3544 470652 3596
rect 483756 3544 483808 3596
rect 498200 3544 498252 3596
rect 511264 3612 511316 3664
rect 513288 3612 513340 3664
rect 575112 3612 575164 3664
rect 514760 3544 514812 3596
rect 517336 3544 517388 3596
rect 582196 3544 582248 3596
rect 4068 3476 4120 3528
rect 1676 3408 1728 3460
rect 11704 3408 11756 3460
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 25504 3476 25556 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 24216 3408 24268 3460
rect 15936 3340 15988 3392
rect 22744 3340 22796 3392
rect 6460 3272 6512 3324
rect 7564 3272 7616 3324
rect 28908 3340 28960 3392
rect 135260 3476 135312 3528
rect 136456 3476 136508 3528
rect 138848 3476 138900 3528
rect 139308 3476 139360 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 402980 3476 403032 3528
rect 408408 3476 408460 3528
rect 135444 3408 135496 3460
rect 139492 3408 139544 3460
rect 142436 3408 142488 3460
rect 143448 3408 143500 3460
rect 145932 3408 145984 3460
rect 403072 3408 403124 3460
rect 404820 3408 404872 3460
rect 461584 3476 461636 3528
rect 462228 3476 462280 3528
rect 465172 3476 465224 3528
rect 466368 3476 466420 3528
rect 468668 3476 468720 3528
rect 469128 3476 469180 3528
rect 472256 3476 472308 3528
rect 473268 3476 473320 3528
rect 479340 3476 479392 3528
rect 480168 3476 480220 3528
rect 486424 3476 486476 3528
rect 487068 3476 487120 3528
rect 501604 3476 501656 3528
rect 469404 3408 469456 3460
rect 471244 3408 471296 3460
rect 502984 3408 503036 3460
rect 504364 3476 504416 3528
rect 505376 3476 505428 3528
rect 507124 3476 507176 3528
rect 508872 3476 508924 3528
rect 514576 3476 514628 3528
rect 578608 3476 578660 3528
rect 510068 3408 510120 3460
rect 514668 3408 514720 3460
rect 579804 3408 579856 3460
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 41880 3340 41932 3392
rect 42984 3340 43036 3392
rect 51356 3340 51408 3392
rect 52368 3340 52420 3392
rect 58440 3340 58492 3392
rect 59268 3340 59320 3392
rect 60832 3340 60884 3392
rect 61936 3340 61988 3392
rect 65524 3340 65576 3392
rect 66168 3340 66220 3392
rect 75000 3340 75052 3392
rect 75828 3340 75880 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 92756 3340 92808 3392
rect 93952 3272 94004 3324
rect 95148 3272 95200 3324
rect 99840 3272 99892 3324
rect 100668 3272 100720 3324
rect 153016 3340 153068 3392
rect 163688 3340 163740 3392
rect 164148 3340 164200 3392
rect 164884 3340 164936 3392
rect 165528 3340 165580 3392
rect 167184 3340 167236 3392
rect 168288 3340 168340 3392
rect 173164 3340 173216 3392
rect 173808 3340 173860 3392
rect 174268 3340 174320 3392
rect 175188 3340 175240 3392
rect 180248 3340 180300 3392
rect 180708 3340 180760 3392
rect 181444 3340 181496 3392
rect 182088 3340 182140 3392
rect 184940 3340 184992 3392
rect 186228 3340 186280 3392
rect 188528 3340 188580 3392
rect 188988 3340 189040 3392
rect 192024 3340 192076 3392
rect 192944 3340 192996 3392
rect 199108 3340 199160 3392
rect 199936 3340 199988 3392
rect 206192 3340 206244 3392
rect 206744 3340 206796 3392
rect 209780 3340 209832 3392
rect 211068 3340 211120 3392
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 245200 3340 245252 3392
rect 246396 3340 246448 3392
rect 258264 3340 258316 3392
rect 259276 3340 259328 3392
rect 262956 3340 263008 3392
rect 264336 3340 264388 3392
rect 276020 3340 276072 3392
rect 277124 3340 277176 3392
rect 280712 3340 280764 3392
rect 281264 3340 281316 3392
rect 291384 3340 291436 3392
rect 292488 3340 292540 3392
rect 298468 3340 298520 3392
rect 300124 3340 300176 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 319720 3340 319772 3392
rect 323584 3340 323636 3392
rect 326804 3340 326856 3392
rect 353944 3340 353996 3392
rect 387156 3340 387208 3392
rect 463792 3340 463844 3392
rect 493968 3340 494020 3392
rect 500592 3340 500644 3392
rect 506388 3340 506440 3392
rect 546684 3340 546736 3392
rect 96252 3204 96304 3256
rect 103336 3204 103388 3256
rect 153292 3272 153344 3324
rect 175464 3272 175516 3324
rect 179512 3272 179564 3324
rect 184204 3272 184256 3324
rect 186136 3272 186188 3324
rect 287796 3272 287848 3324
rect 294604 3272 294656 3324
rect 337476 3272 337528 3324
rect 345664 3272 345716 3324
rect 348056 3272 348108 3324
rect 374644 3272 374696 3324
rect 390652 3272 390704 3324
rect 465264 3272 465316 3324
rect 505008 3272 505060 3324
rect 543188 3272 543240 3324
rect 106924 3136 106976 3188
rect 153200 3204 153252 3256
rect 171968 3204 172020 3256
rect 177304 3204 177356 3256
rect 394240 3204 394292 3256
rect 466644 3204 466696 3256
rect 503628 3204 503680 3256
rect 539600 3204 539652 3256
rect 12348 3068 12400 3120
rect 14464 3068 14516 3120
rect 30104 3068 30156 3120
rect 32404 3068 32456 3120
rect 110512 3068 110564 3120
rect 155960 3136 156012 3188
rect 183744 3136 183796 3188
rect 188344 3136 188396 3188
rect 284300 3136 284352 3188
rect 285588 3136 285640 3188
rect 316224 3136 316276 3188
rect 322296 3136 322348 3188
rect 397736 3136 397788 3188
rect 466552 3136 466604 3188
rect 493876 3136 493928 3188
rect 497096 3136 497148 3188
rect 503536 3136 503588 3188
rect 536104 3136 536156 3188
rect 67916 3000 67968 3052
rect 71228 3000 71280 3052
rect 114008 3000 114060 3052
rect 156052 3068 156104 3120
rect 176660 3068 176712 3120
rect 180064 3068 180116 3120
rect 231032 3068 231084 3120
rect 233884 3068 233936 3120
rect 426164 3068 426216 3120
rect 474832 3068 474884 3120
rect 485044 3068 485096 3120
rect 487620 3068 487672 3120
rect 502248 3068 502300 3120
rect 532516 3068 532568 3120
rect 117596 2932 117648 2984
rect 157432 3000 157484 3052
rect 248788 3000 248840 3052
rect 251824 3000 251876 3052
rect 415492 3000 415544 3052
rect 121092 2864 121144 2916
rect 157340 2932 157392 2984
rect 223948 2932 224000 2984
rect 224776 2932 224828 2984
rect 433248 2932 433300 2984
rect 476304 3000 476356 3052
rect 497464 3000 497516 3052
rect 499396 3000 499448 3052
rect 500868 3000 500920 3052
rect 529020 3000 529072 3052
rect 447416 2932 447468 2984
rect 448428 2932 448480 2984
rect 158812 2864 158864 2916
rect 436744 2864 436796 2916
rect 476212 2932 476264 2984
rect 490564 2932 490616 2984
rect 492312 2932 492364 2984
rect 500776 2932 500828 2984
rect 525432 2932 525484 2984
rect 124680 2796 124732 2848
rect 160192 2796 160244 2848
rect 440332 2796 440384 2848
rect 441528 2796 441580 2848
rect 443828 2796 443880 2848
rect 478972 2864 479024 2916
rect 499488 2864 499540 2916
rect 521844 2864 521896 2916
rect 450912 2796 450964 2848
rect 480260 2796 480312 2848
rect 499304 2796 499356 2848
rect 518348 2796 518400 2848
rect 340880 1912 340932 1964
rect 342168 1912 342220 1964
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 637566 3464 697303
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 637560 3476 637566
rect 3424 637502 3476 637508
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3436 583710 3464 632023
rect 3528 626550 3556 684247
rect 3606 671256 3662 671265
rect 3606 671191 3662 671200
rect 3516 626544 3568 626550
rect 3516 626486 3568 626492
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 583704 3476 583710
rect 3424 583646 3476 583652
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 539578 3464 579935
rect 3528 572694 3556 619103
rect 3620 615466 3648 671191
rect 3698 658200 3754 658209
rect 3698 658135 3754 658144
rect 3608 615460 3660 615466
rect 3608 615402 3660 615408
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3516 572688 3568 572694
rect 3516 572630 3568 572636
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 539572 3476 539578
rect 3424 539514 3476 539520
rect 3528 528562 3556 566879
rect 3620 561678 3648 606047
rect 3712 605810 3740 658135
rect 3790 645144 3846 645153
rect 3790 645079 3846 645088
rect 3700 605804 3752 605810
rect 3700 605746 3752 605752
rect 3804 594794 3832 645079
rect 8220 642394 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 642462 24808 699654
rect 41340 642530 41368 700334
rect 56796 700194 56824 703520
rect 72988 702434 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72988 702406 73108 702434
rect 56784 700188 56836 700194
rect 56784 700130 56836 700136
rect 57888 700188 57940 700194
rect 57888 700130 57940 700136
rect 57900 642598 57928 700130
rect 57888 642592 57940 642598
rect 57888 642534 57940 642540
rect 41328 642524 41380 642530
rect 41328 642466 41380 642472
rect 24768 642456 24820 642462
rect 24768 642398 24820 642404
rect 73080 642394 73108 702406
rect 89640 642462 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 106200 642530 106228 700334
rect 121656 699718 121684 703520
rect 137848 702434 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137848 702406 137968 702434
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 122760 642598 122788 699654
rect 110144 642592 110196 642598
rect 110144 642534 110196 642540
rect 122748 642592 122800 642598
rect 122748 642534 122800 642540
rect 97356 642524 97408 642530
rect 97356 642466 97408 642472
rect 106188 642524 106240 642530
rect 106188 642466 106240 642472
rect 84660 642456 84712 642462
rect 84660 642398 84712 642404
rect 89628 642456 89680 642462
rect 89628 642398 89680 642404
rect 8208 642388 8260 642394
rect 8208 642330 8260 642336
rect 72792 642388 72844 642394
rect 72792 642330 72844 642336
rect 73068 642388 73120 642394
rect 73068 642330 73120 642336
rect 72804 639282 72832 642330
rect 84672 639282 84700 642398
rect 97368 639282 97396 642466
rect 110156 639282 110184 642534
rect 135536 642456 135588 642462
rect 135536 642398 135588 642404
rect 122840 642388 122892 642394
rect 122840 642330 122892 642336
rect 122852 639282 122880 642330
rect 72804 639254 72874 639282
rect 84672 639254 84734 639282
rect 97368 639254 97434 639282
rect 72846 638996 72874 639254
rect 84706 638996 84734 639254
rect 97406 638996 97434 639254
rect 110126 639254 110184 639282
rect 122846 639254 122880 639282
rect 135548 639282 135576 642398
rect 137940 642394 137968 702406
rect 148232 642524 148284 642530
rect 148232 642466 148284 642472
rect 137928 642388 137980 642394
rect 137928 642330 137980 642336
rect 148244 639282 148272 642466
rect 154500 642462 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 161020 642592 161072 642598
rect 161020 642534 161072 642540
rect 154488 642456 154540 642462
rect 154488 642398 154540 642404
rect 161032 639282 161060 642534
rect 171060 642530 171088 700198
rect 186516 700194 186544 703520
rect 186504 700188 186556 700194
rect 186504 700130 186556 700136
rect 187608 700188 187660 700194
rect 187608 700130 187660 700136
rect 171048 642524 171100 642530
rect 171048 642466 171100 642472
rect 186412 642456 186464 642462
rect 186412 642398 186464 642404
rect 173716 642388 173768 642394
rect 173716 642330 173768 642336
rect 173728 639282 173756 642330
rect 135548 639254 135594 639282
rect 148244 639254 148314 639282
rect 110126 638996 110154 639254
rect 122846 638996 122874 639254
rect 135566 638996 135594 639254
rect 148286 638996 148314 639254
rect 161006 639254 161060 639282
rect 173726 639254 173756 639282
rect 186424 639282 186452 642398
rect 187620 642394 187648 700130
rect 199108 642524 199160 642530
rect 199108 642466 199160 642472
rect 187608 642388 187660 642394
rect 187608 642330 187660 642336
rect 199120 639282 199148 642466
rect 202800 642462 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 642456 202840 642462
rect 202788 642398 202840 642404
rect 219360 642394 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 235920 642462 235948 700334
rect 251468 700126 251496 703520
rect 251456 700120 251508 700126
rect 251456 700062 251508 700068
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 224592 642456 224644 642462
rect 224592 642398 224644 642404
rect 235908 642456 235960 642462
rect 235908 642398 235960 642404
rect 249984 642456 250036 642462
rect 249984 642398 250036 642404
rect 211896 642388 211948 642394
rect 211896 642330 211948 642336
rect 219348 642388 219400 642394
rect 219348 642330 219400 642336
rect 211908 639282 211936 642330
rect 186424 639254 186474 639282
rect 199120 639254 199194 639282
rect 161006 638996 161034 639254
rect 173726 638996 173754 639254
rect 186446 638996 186474 639254
rect 199166 638996 199194 639254
rect 211886 639254 211936 639282
rect 224604 639282 224632 642398
rect 237288 642388 237340 642394
rect 237288 642330 237340 642336
rect 237300 639282 237328 642330
rect 249996 639282 250024 642398
rect 252480 642394 252508 700062
rect 267660 642394 267688 703520
rect 283852 700126 283880 703520
rect 283840 700120 283892 700126
rect 283840 700062 283892 700068
rect 284944 700120 284996 700126
rect 284944 700062 284996 700068
rect 284956 643074 284984 700062
rect 300136 699718 300164 703520
rect 316328 699718 316356 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 364996 700330 365024 703520
rect 378048 700392 378100 700398
rect 378048 700334 378100 700340
rect 339408 700324 339460 700330
rect 339408 700266 339460 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 351828 700324 351880 700330
rect 351828 700266 351880 700272
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 365628 700324 365680 700330
rect 365628 700266 365680 700272
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 314568 699712 314620 699718
rect 314568 699654 314620 699660
rect 316316 699712 316368 699718
rect 316316 699654 316368 699660
rect 327724 699712 327776 699718
rect 327724 699654 327776 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 284944 643068 284996 643074
rect 284944 643010 284996 643016
rect 288164 643068 288216 643074
rect 288164 643010 288216 643016
rect 252468 642388 252520 642394
rect 252468 642330 252520 642336
rect 262772 642388 262824 642394
rect 262772 642330 262824 642336
rect 267648 642388 267700 642394
rect 267648 642330 267700 642336
rect 275468 642388 275520 642394
rect 275468 642330 275520 642336
rect 262784 639282 262812 642330
rect 224604 639254 224634 639282
rect 237300 639254 237354 639282
rect 249996 639254 250074 639282
rect 211886 638996 211914 639254
rect 224606 638996 224634 639254
rect 237326 638996 237354 639254
rect 250046 638996 250074 639254
rect 262766 639254 262812 639282
rect 275480 639282 275508 642330
rect 288176 639282 288204 643010
rect 300780 641730 300808 699654
rect 314580 641782 314608 699654
rect 327736 641782 327764 699654
rect 313648 641776 313700 641782
rect 300780 641702 300900 641730
rect 313648 641718 313700 641724
rect 314568 641776 314620 641782
rect 314568 641718 314620 641724
rect 326344 641776 326396 641782
rect 326344 641718 326396 641724
rect 327724 641776 327776 641782
rect 327724 641718 327776 641724
rect 300872 639282 300900 641702
rect 313660 639282 313688 641718
rect 275480 639254 275514 639282
rect 288176 639254 288234 639282
rect 300872 639254 300954 639282
rect 262766 638996 262794 639254
rect 275486 638996 275514 639254
rect 288206 638996 288234 639254
rect 300926 638996 300954 639254
rect 313646 639254 313688 639282
rect 326356 639282 326384 641718
rect 339420 639282 339448 700266
rect 351840 639282 351868 700266
rect 365640 641782 365668 700266
rect 378060 641782 378088 700334
rect 381188 700330 381216 703520
rect 397472 700398 397500 703520
rect 402888 700460 402940 700466
rect 402888 700402 402940 700408
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 381176 700324 381228 700330
rect 381176 700266 381228 700272
rect 390468 700324 390520 700330
rect 390468 700266 390520 700272
rect 390480 641782 390508 700266
rect 364524 641776 364576 641782
rect 364524 641718 364576 641724
rect 365628 641776 365680 641782
rect 365628 641718 365680 641724
rect 377220 641776 377272 641782
rect 377220 641718 377272 641724
rect 378048 641776 378100 641782
rect 378048 641718 378100 641724
rect 390008 641776 390060 641782
rect 390008 641718 390060 641724
rect 390468 641776 390520 641782
rect 390468 641718 390520 641724
rect 364536 639282 364564 641718
rect 326356 639254 326394 639282
rect 313646 638996 313674 639254
rect 326366 638996 326394 639254
rect 339086 639254 339448 639282
rect 351806 639254 351868 639282
rect 364526 639254 364564 639282
rect 377232 639282 377260 641718
rect 390020 639282 390048 641718
rect 402900 639282 402928 700402
rect 413664 700330 413692 703520
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 441528 700460 441580 700466
rect 441528 700402 441580 700408
rect 416688 700392 416740 700398
rect 416688 700334 416740 700340
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 416700 641782 416728 700334
rect 429108 700324 429160 700330
rect 429108 700266 429160 700272
rect 429120 641782 429148 700266
rect 441540 642598 441568 700402
rect 446140 700398 446168 703520
rect 446128 700392 446180 700398
rect 446128 700334 446180 700340
rect 453948 700392 454000 700398
rect 453948 700334 454000 700340
rect 440884 642592 440936 642598
rect 440884 642534 440936 642540
rect 441528 642592 441580 642598
rect 441528 642534 441580 642540
rect 415400 641776 415452 641782
rect 415400 641718 415452 641724
rect 416688 641776 416740 641782
rect 416688 641718 416740 641724
rect 428096 641776 428148 641782
rect 428096 641718 428148 641724
rect 429108 641776 429160 641782
rect 429108 641718 429160 641724
rect 415412 639282 415440 641718
rect 377232 639254 377274 639282
rect 339086 638996 339114 639254
rect 351806 638996 351834 639254
rect 364526 638996 364554 639254
rect 377246 638996 377274 639254
rect 389966 639254 390048 639282
rect 402686 639254 402928 639282
rect 415406 639254 415440 639282
rect 428108 639282 428136 641718
rect 440896 639282 440924 642534
rect 453960 639282 453988 700334
rect 462332 700330 462360 703520
rect 478524 700466 478552 703520
rect 480168 700528 480220 700534
rect 480168 700470 480220 700476
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 466368 700324 466420 700330
rect 466368 700266 466420 700272
rect 466380 639282 466408 700266
rect 480180 641782 480208 700470
rect 492588 700460 492640 700466
rect 492588 700402 492640 700408
rect 492600 641782 492628 700402
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 505008 700392 505060 700398
rect 505008 700334 505060 700340
rect 505020 641782 505048 700334
rect 511000 700330 511028 703520
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 575860 700330 575888 703520
rect 510988 700324 511040 700330
rect 510988 700266 511040 700272
rect 517428 700324 517480 700330
rect 517428 700266 517480 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 517440 641782 517468 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 519544 696992 519596 696998
rect 519544 696934 519596 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 478972 641776 479024 641782
rect 478972 641718 479024 641724
rect 480168 641776 480220 641782
rect 480168 641718 480220 641724
rect 491760 641776 491812 641782
rect 491760 641718 491812 641724
rect 492588 641776 492640 641782
rect 492588 641718 492640 641724
rect 504456 641776 504508 641782
rect 504456 641718 504508 641724
rect 505008 641776 505060 641782
rect 505008 641718 505060 641724
rect 516508 641776 516560 641782
rect 516508 641718 516560 641724
rect 517428 641776 517480 641782
rect 517428 641718 517480 641724
rect 428108 639254 428154 639282
rect 389966 638996 389994 639254
rect 402686 638996 402714 639254
rect 415406 638996 415434 639254
rect 428126 638996 428154 639254
rect 440846 639254 440924 639282
rect 453566 639254 453988 639282
rect 466286 639254 466408 639282
rect 478984 639282 479012 641718
rect 491772 639282 491800 641718
rect 504468 639282 504496 641718
rect 516520 639282 516548 641718
rect 478984 639254 479034 639282
rect 440846 638996 440874 639254
rect 453566 638996 453594 639254
rect 466286 638996 466314 639254
rect 479006 638996 479034 639254
rect 491726 639254 491800 639282
rect 504446 639254 504496 639282
rect 516466 639254 516548 639282
rect 491726 638996 491754 639254
rect 504446 638996 504474 639254
rect 516466 638996 516494 639254
rect 69020 637560 69072 637566
rect 69020 637502 69072 637508
rect 69032 636721 69060 637502
rect 519556 636857 519584 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 519636 683188 519688 683194
rect 519636 683130 519688 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 519542 636848 519598 636857
rect 519542 636783 519598 636792
rect 69018 636712 69074 636721
rect 69018 636647 69074 636656
rect 519544 630692 519596 630698
rect 519544 630634 519596 630640
rect 69020 626544 69072 626550
rect 69020 626486 69072 626492
rect 69032 626385 69060 626486
rect 69018 626376 69074 626385
rect 69018 626311 69074 626320
rect 69018 615496 69074 615505
rect 69018 615431 69020 615440
rect 69072 615431 69074 615440
rect 69020 615402 69072 615408
rect 69020 605804 69072 605810
rect 69020 605746 69072 605752
rect 69032 604625 69060 605746
rect 69018 604616 69074 604625
rect 69018 604551 69074 604560
rect 3792 594788 3844 594794
rect 3792 594730 3844 594736
rect 69020 594788 69072 594794
rect 69020 594730 69072 594736
rect 69032 593745 69060 594730
rect 69018 593736 69074 593745
rect 69018 593671 69074 593680
rect 3698 593056 3754 593065
rect 3698 592991 3754 593000
rect 3608 561672 3660 561678
rect 3608 561614 3660 561620
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3516 528556 3568 528562
rect 3516 528498 3568 528504
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 496806 3464 527847
rect 3620 517478 3648 553823
rect 3712 550594 3740 592991
rect 69020 583704 69072 583710
rect 69020 583646 69072 583652
rect 69032 582865 69060 583646
rect 69018 582856 69074 582865
rect 69018 582791 69074 582800
rect 519556 581777 519584 630634
rect 519648 626249 519676 683130
rect 519728 670744 519780 670750
rect 580172 670744 580224 670750
rect 519728 670686 519780 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 519634 626240 519690 626249
rect 519634 626175 519690 626184
rect 519636 616888 519688 616894
rect 519636 616830 519688 616836
rect 519542 581768 519598 581777
rect 519542 581703 519598 581712
rect 519544 576904 519596 576910
rect 519544 576846 519596 576852
rect 69020 572688 69072 572694
rect 69020 572630 69072 572636
rect 69032 571985 69060 572630
rect 69018 571976 69074 571985
rect 69018 571911 69074 571920
rect 69020 561672 69072 561678
rect 69020 561614 69072 561620
rect 69032 560969 69060 561614
rect 69018 560960 69074 560969
rect 69018 560895 69074 560904
rect 3700 550588 3752 550594
rect 3700 550530 3752 550536
rect 69020 550588 69072 550594
rect 69020 550530 69072 550536
rect 69032 550225 69060 550530
rect 69018 550216 69074 550225
rect 69018 550151 69074 550160
rect 3698 540832 3754 540841
rect 3698 540767 3754 540776
rect 3608 517472 3660 517478
rect 3608 517414 3660 517420
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 496800 3476 496806
rect 3424 496742 3476 496748
rect 3422 488744 3478 488753
rect 3422 488679 3478 488688
rect 3436 463690 3464 488679
rect 3528 485790 3556 514791
rect 3712 507822 3740 540767
rect 69020 539572 69072 539578
rect 69020 539514 69072 539520
rect 69032 539209 69060 539514
rect 69018 539200 69074 539209
rect 69018 539135 69074 539144
rect 519556 537441 519584 576846
rect 519648 570625 519676 616830
rect 519740 615097 519768 670686
rect 580170 670647 580226 670656
rect 580170 657384 580226 657393
rect 580170 657319 580226 657328
rect 580184 656946 580212 657319
rect 519820 656940 519872 656946
rect 519820 656882 519872 656888
rect 580172 656940 580224 656946
rect 580172 656882 580224 656888
rect 519726 615088 519782 615097
rect 519726 615023 519782 615032
rect 519832 603945 519860 656882
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 519912 643136 519964 643142
rect 519912 643078 519964 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 519818 603936 519874 603945
rect 519818 603871 519874 603880
rect 519728 603152 519780 603158
rect 519728 603094 519780 603100
rect 519634 570616 519690 570625
rect 519634 570551 519690 570560
rect 519636 563100 519688 563106
rect 519636 563042 519688 563048
rect 519542 537432 519598 537441
rect 519542 537367 519598 537376
rect 69020 528556 69072 528562
rect 69020 528498 69072 528504
rect 69032 528329 69060 528498
rect 69018 528320 69074 528329
rect 69018 528255 69074 528264
rect 519648 526289 519676 563042
rect 519740 559609 519768 603094
rect 519924 592929 519952 643078
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 519910 592920 519966 592929
rect 519910 592855 519966 592864
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 519820 590708 519872 590714
rect 519820 590650 519872 590656
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 519726 559600 519782 559609
rect 519726 559535 519782 559544
rect 519728 550656 519780 550662
rect 519728 550598 519780 550604
rect 519634 526280 519690 526289
rect 519634 526215 519690 526224
rect 519544 524476 519596 524482
rect 519544 524418 519596 524424
rect 69020 517472 69072 517478
rect 69018 517440 69020 517449
rect 69072 517440 69074 517449
rect 69018 517375 69074 517384
rect 3700 507816 3752 507822
rect 3700 507758 3752 507764
rect 69020 507816 69072 507822
rect 69020 507758 69072 507764
rect 69032 506569 69060 507758
rect 69018 506560 69074 506569
rect 69018 506495 69074 506504
rect 3606 501800 3662 501809
rect 3606 501735 3662 501744
rect 3516 485784 3568 485790
rect 3516 485726 3568 485732
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3424 463684 3476 463690
rect 3424 463626 3476 463632
rect 3528 452606 3556 475623
rect 3620 474706 3648 501735
rect 69020 496800 69072 496806
rect 69020 496742 69072 496748
rect 69032 495689 69060 496742
rect 69018 495680 69074 495689
rect 69018 495615 69074 495624
rect 519556 492833 519584 524418
rect 519740 515137 519768 550598
rect 519832 548457 519860 590650
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 551168 580226 551177
rect 580170 551103 580226 551112
rect 580184 550662 580212 551103
rect 580172 550656 580224 550662
rect 580172 550598 580224 550604
rect 519818 548448 519874 548457
rect 519818 548383 519874 548392
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 519820 536852 519872 536858
rect 519820 536794 519872 536800
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 519726 515128 519782 515137
rect 519726 515063 519782 515072
rect 519636 510672 519688 510678
rect 519636 510614 519688 510620
rect 519542 492824 519598 492833
rect 519542 492759 519598 492768
rect 69020 485784 69072 485790
rect 69020 485726 69072 485732
rect 69032 484809 69060 485726
rect 69018 484800 69074 484809
rect 69018 484735 69074 484744
rect 519544 484424 519596 484430
rect 519544 484366 519596 484372
rect 3608 474700 3660 474706
rect 3608 474642 3660 474648
rect 69020 474700 69072 474706
rect 69020 474642 69072 474648
rect 69032 473929 69060 474642
rect 69018 473920 69074 473929
rect 69018 473855 69074 473864
rect 69020 463684 69072 463690
rect 69020 463626 69072 463632
rect 69032 463049 69060 463626
rect 69018 463040 69074 463049
rect 69018 462975 69074 462984
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3516 452600 3568 452606
rect 3516 452542 3568 452548
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3436 430574 3464 449511
rect 3620 441590 3648 462567
rect 519556 459649 519584 484366
rect 519648 481817 519676 510614
rect 519832 504121 519860 536794
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 519818 504112 519874 504121
rect 519818 504047 519874 504056
rect 580170 497992 580226 498001
rect 580170 497927 580226 497936
rect 580184 496874 580212 497927
rect 519728 496868 519780 496874
rect 519728 496810 519780 496816
rect 580172 496868 580224 496874
rect 580172 496810 580224 496816
rect 519634 481808 519690 481817
rect 519634 481743 519690 481752
rect 519740 470801 519768 496810
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 519726 470792 519782 470801
rect 519726 470727 519782 470736
rect 580000 470626 580028 471407
rect 519636 470620 519688 470626
rect 519636 470562 519688 470568
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 519542 459640 519598 459649
rect 519542 459575 519598 459584
rect 519544 456816 519596 456822
rect 519544 456758 519596 456764
rect 69020 452600 69072 452606
rect 69020 452542 69072 452548
rect 69032 452169 69060 452542
rect 69018 452160 69074 452169
rect 69018 452095 69074 452104
rect 3608 441584 3660 441590
rect 3608 441526 3660 441532
rect 69020 441584 69072 441590
rect 69020 441526 69072 441532
rect 69032 441289 69060 441526
rect 69018 441280 69074 441289
rect 69018 441215 69074 441224
rect 519556 437481 519584 456758
rect 519648 448633 519676 470562
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 519634 448624 519690 448633
rect 519634 448559 519690 448568
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 519636 444440 519688 444446
rect 519636 444382 519688 444388
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 519542 437472 519598 437481
rect 519542 437407 519598 437416
rect 3514 436656 3570 436665
rect 3514 436591 3570 436600
rect 3424 430568 3476 430574
rect 3424 430510 3476 430516
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 409834 3464 423535
rect 3528 419490 3556 436591
rect 519544 430636 519596 430642
rect 519544 430578 519596 430584
rect 69020 430568 69072 430574
rect 69020 430510 69072 430516
rect 69032 430409 69060 430510
rect 69018 430400 69074 430409
rect 69018 430335 69074 430344
rect 3516 419484 3568 419490
rect 3516 419426 3568 419432
rect 69020 419484 69072 419490
rect 69020 419426 69072 419432
rect 69032 419393 69060 419426
rect 69018 419384 69074 419393
rect 69018 419319 69074 419328
rect 519556 415313 519584 430578
rect 519648 426329 519676 444382
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 519634 426320 519690 426329
rect 519634 426255 519690 426264
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 519636 418192 519688 418198
rect 519636 418134 519688 418140
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 519542 415304 519598 415313
rect 519542 415239 519598 415248
rect 3514 410544 3570 410553
rect 3514 410479 3570 410488
rect 3424 409828 3476 409834
rect 3424 409770 3476 409776
rect 3528 398818 3556 410479
rect 69020 409828 69072 409834
rect 69020 409770 69072 409776
rect 69032 408649 69060 409770
rect 69018 408640 69074 408649
rect 69018 408575 69074 408584
rect 519544 404388 519596 404394
rect 519544 404330 519596 404336
rect 3516 398812 3568 398818
rect 3516 398754 3568 398760
rect 69020 398812 69072 398818
rect 69020 398754 69072 398760
rect 69032 397633 69060 398754
rect 69018 397624 69074 397633
rect 69018 397559 69074 397568
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 387802 3464 397423
rect 519556 393009 519584 404330
rect 519648 404161 519676 418134
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 519634 404152 519690 404161
rect 519634 404087 519690 404096
rect 519542 393000 519598 393009
rect 519542 392935 519598 392944
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 580184 390590 580212 391711
rect 519544 390584 519596 390590
rect 519544 390526 519596 390532
rect 580172 390584 580224 390590
rect 580172 390526 580224 390532
rect 3424 387796 3476 387802
rect 3424 387738 3476 387744
rect 69020 387796 69072 387802
rect 69020 387738 69072 387744
rect 69032 386753 69060 387738
rect 69018 386744 69074 386753
rect 69018 386679 69074 386688
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 376718 3464 384367
rect 519556 381993 519584 390526
rect 519542 381984 519598 381993
rect 519542 381919 519598 381928
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 519544 378208 519596 378214
rect 519544 378150 519596 378156
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 3424 376712 3476 376718
rect 3424 376654 3476 376660
rect 69020 376712 69072 376718
rect 69020 376654 69072 376660
rect 69032 375873 69060 376654
rect 69018 375864 69074 375873
rect 69018 375799 69074 375808
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 365702 3464 371311
rect 519556 370841 519584 378150
rect 519542 370832 519598 370841
rect 519542 370767 519598 370776
rect 3424 365696 3476 365702
rect 3424 365638 3476 365644
rect 69020 365696 69072 365702
rect 69020 365638 69072 365644
rect 69032 364993 69060 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 69018 364984 69074 364993
rect 69018 364919 69074 364928
rect 580184 364410 580212 365055
rect 519360 364404 519412 364410
rect 519360 364346 519412 364352
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 519372 359825 519400 364346
rect 519358 359816 519414 359825
rect 519358 359751 519414 359760
rect 3422 358456 3478 358465
rect 3422 358391 3478 358400
rect 3436 354686 3464 358391
rect 3424 354680 3476 354686
rect 3424 354622 3476 354628
rect 69020 354680 69072 354686
rect 69020 354622 69072 354628
rect 69032 354113 69060 354622
rect 69018 354104 69074 354113
rect 69018 354039 69074 354048
rect 519820 351960 519872 351966
rect 580172 351960 580224 351966
rect 519820 351902 519872 351908
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 519832 348673 519860 351902
rect 580170 351863 580226 351872
rect 519818 348664 519874 348673
rect 519818 348599 519874 348608
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3160 343602 3188 345335
rect 3148 343596 3200 343602
rect 3148 343538 3200 343544
rect 69020 343596 69072 343602
rect 69020 343538 69072 343544
rect 69032 343233 69060 343538
rect 69018 343224 69074 343233
rect 69018 343159 69074 343168
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 580184 338162 580212 338535
rect 520004 338156 520056 338162
rect 520004 338098 520056 338104
rect 580172 338156 580224 338162
rect 580172 338098 580224 338104
rect 520016 337521 520044 338098
rect 520002 337512 520058 337521
rect 520002 337447 520058 337456
rect 3422 332344 3478 332353
rect 3422 332279 3478 332288
rect 3436 331906 3464 332279
rect 69018 332208 69074 332217
rect 69018 332143 69074 332152
rect 69032 331906 69060 332143
rect 3424 331900 3476 331906
rect 3424 331842 3476 331848
rect 69020 331900 69072 331906
rect 69020 331842 69072 331848
rect 519358 326360 519414 326369
rect 519358 326295 519414 326304
rect 519372 325650 519400 326295
rect 519360 325644 519412 325650
rect 519360 325586 519412 325592
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 69018 321328 69074 321337
rect 69018 321263 69074 321272
rect 69032 320210 69060 321263
rect 3424 320204 3476 320210
rect 3424 320146 3476 320152
rect 69020 320204 69072 320210
rect 69020 320146 69072 320152
rect 3436 319297 3464 320146
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 520186 315344 520242 315353
rect 520186 315279 520242 315288
rect 520200 313274 520228 315279
rect 520188 313268 520240 313274
rect 520188 313210 520240 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 69018 310448 69074 310457
rect 69018 310383 69074 310392
rect 69032 309194 69060 310383
rect 3424 309188 3476 309194
rect 3424 309130 3476 309136
rect 69020 309188 69072 309194
rect 69020 309130 69072 309136
rect 3436 306241 3464 309130
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 519358 304192 519414 304201
rect 519358 304127 519414 304136
rect 69018 299568 69074 299577
rect 3424 299532 3476 299538
rect 69018 299503 69020 299512
rect 3424 299474 3476 299480
rect 69072 299503 69074 299512
rect 69020 299474 69072 299480
rect 3436 293185 3464 299474
rect 519372 299470 519400 304127
rect 519360 299464 519412 299470
rect 519360 299406 519412 299412
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 519542 293176 519598 293185
rect 519542 293111 519598 293120
rect 69018 288688 69074 288697
rect 69018 288623 69074 288632
rect 69032 288454 69060 288623
rect 3424 288448 3476 288454
rect 3424 288390 3476 288396
rect 69020 288448 69072 288454
rect 69020 288390 69072 288396
rect 3436 280129 3464 288390
rect 519556 285666 519584 293111
rect 519544 285660 519596 285666
rect 519544 285602 519596 285608
rect 580172 285660 580224 285666
rect 580172 285602 580224 285608
rect 580184 285433 580212 285602
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 519542 282024 519598 282033
rect 519542 281959 519598 281968
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 69018 277808 69074 277817
rect 69018 277743 69074 277752
rect 69032 277438 69060 277743
rect 3516 277432 3568 277438
rect 3516 277374 3568 277380
rect 69020 277432 69072 277438
rect 69020 277374 69072 277380
rect 3528 267209 3556 277374
rect 519556 273222 519584 281959
rect 519544 273216 519596 273222
rect 519544 273158 519596 273164
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 519542 270872 519598 270881
rect 519542 270807 519598 270816
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 69018 266928 69074 266937
rect 69018 266863 69074 266872
rect 69032 266422 69060 266863
rect 3424 266416 3476 266422
rect 3424 266358 3476 266364
rect 69020 266416 69072 266422
rect 69020 266358 69072 266364
rect 3436 254153 3464 266358
rect 519556 259418 519584 270807
rect 519634 259856 519690 259865
rect 519634 259791 519690 259800
rect 519544 259412 519596 259418
rect 519544 259354 519596 259360
rect 69018 256048 69074 256057
rect 69018 255983 69074 255992
rect 69032 255338 69060 255983
rect 3516 255332 3568 255338
rect 3516 255274 3568 255280
rect 69020 255332 69072 255338
rect 69020 255274 69072 255280
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 244316 3476 244322
rect 3424 244258 3476 244264
rect 3436 228041 3464 244258
rect 3528 241097 3556 255274
rect 519542 248704 519598 248713
rect 519542 248639 519598 248648
rect 69018 245168 69074 245177
rect 69018 245103 69074 245112
rect 69032 244322 69060 245103
rect 69020 244316 69072 244322
rect 69020 244258 69072 244264
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 69018 234288 69074 234297
rect 69018 234223 69074 234232
rect 69032 233306 69060 234223
rect 3516 233300 3568 233306
rect 3516 233242 3568 233248
rect 69020 233300 69072 233306
rect 69020 233242 69072 233248
rect 3422 228032 3478 228041
rect 3422 227967 3478 227976
rect 3424 222216 3476 222222
rect 3424 222158 3476 222164
rect 3436 201929 3464 222158
rect 3528 214985 3556 233242
rect 519556 233238 519584 248639
rect 519648 245614 519676 259791
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 519636 245608 519688 245614
rect 580172 245608 580224 245614
rect 519636 245550 519688 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 519634 237552 519690 237561
rect 519634 237487 519690 237496
rect 519544 233232 519596 233238
rect 519544 233174 519596 233180
rect 519542 226536 519598 226545
rect 519542 226471 519598 226480
rect 69018 223408 69074 223417
rect 69018 223343 69074 223352
rect 69032 222222 69060 223343
rect 69020 222216 69072 222222
rect 69020 222158 69072 222164
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 69018 212528 69074 212537
rect 69018 212463 69074 212472
rect 69032 211206 69060 212463
rect 3608 211200 3660 211206
rect 3608 211142 3660 211148
rect 69020 211200 69072 211206
rect 69020 211142 69072 211148
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3516 201544 3568 201550
rect 3516 201486 3568 201492
rect 3424 190528 3476 190534
rect 3424 190470 3476 190476
rect 3436 162897 3464 190470
rect 3528 175953 3556 201486
rect 3620 188873 3648 211142
rect 519556 206990 519584 226471
rect 519648 219434 519676 237487
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 519636 219428 519688 219434
rect 519636 219370 519688 219376
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 519726 215384 519782 215393
rect 519726 215319 519782 215328
rect 519544 206984 519596 206990
rect 519544 206926 519596 206932
rect 519634 204368 519690 204377
rect 519634 204303 519690 204312
rect 69018 201648 69074 201657
rect 69018 201583 69074 201592
rect 69032 201550 69060 201583
rect 69020 201544 69072 201550
rect 69020 201486 69072 201492
rect 519542 193216 519598 193225
rect 519542 193151 519598 193160
rect 69018 190632 69074 190641
rect 69018 190567 69074 190576
rect 69032 190534 69060 190567
rect 69020 190528 69072 190534
rect 69020 190470 69072 190476
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 69018 179752 69074 179761
rect 69018 179687 69074 179696
rect 69032 179450 69060 179687
rect 3608 179444 3660 179450
rect 3608 179386 3660 179392
rect 69020 179444 69072 179450
rect 69020 179386 69072 179392
rect 3514 175944 3570 175953
rect 3514 175879 3570 175888
rect 3516 168428 3568 168434
rect 3516 168370 3568 168376
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3424 157412 3476 157418
rect 3424 157354 3476 157360
rect 3436 123729 3464 157354
rect 3528 136785 3556 168370
rect 3620 149841 3648 179386
rect 69018 168872 69074 168881
rect 69018 168807 69074 168816
rect 69032 168434 69060 168807
rect 69020 168428 69072 168434
rect 69020 168370 69072 168376
rect 519556 167006 519584 193151
rect 519648 179382 519676 204303
rect 519740 193186 519768 215319
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 519728 193180 519780 193186
rect 519728 193122 519780 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 519726 182064 519782 182073
rect 519726 181999 519782 182008
rect 519636 179376 519688 179382
rect 519636 179318 519688 179324
rect 519634 171048 519690 171057
rect 519634 170983 519690 170992
rect 519544 167000 519596 167006
rect 519544 166942 519596 166948
rect 519542 159896 519598 159905
rect 519542 159831 519598 159840
rect 69018 157992 69074 158001
rect 69018 157927 69074 157936
rect 69032 157418 69060 157927
rect 69020 157412 69072 157418
rect 69020 157354 69072 157360
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 69018 147112 69074 147121
rect 69018 147047 69074 147056
rect 69032 146334 69060 147047
rect 3700 146328 3752 146334
rect 3700 146270 3752 146276
rect 69020 146328 69072 146334
rect 69020 146270 69072 146276
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3608 135312 3660 135318
rect 3608 135254 3660 135260
rect 3516 124228 3568 124234
rect 3516 124170 3568 124176
rect 3422 123720 3478 123729
rect 3422 123655 3478 123664
rect 3424 113212 3476 113218
rect 3424 113154 3476 113160
rect 3436 71641 3464 113154
rect 3528 84697 3556 124170
rect 3620 97617 3648 135254
rect 3712 110673 3740 146270
rect 69018 136232 69074 136241
rect 69018 136167 69074 136176
rect 69032 135318 69060 136167
rect 69020 135312 69072 135318
rect 69020 135254 69072 135260
rect 519556 126954 519584 159831
rect 519648 139398 519676 170983
rect 519740 153202 519768 181999
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 519728 153196 519780 153202
rect 519728 153138 519780 153144
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 519818 148744 519874 148753
rect 519818 148679 519874 148688
rect 519636 139392 519688 139398
rect 519636 139334 519688 139340
rect 519726 137728 519782 137737
rect 519726 137663 519782 137672
rect 519544 126948 519596 126954
rect 519544 126890 519596 126896
rect 519634 126576 519690 126585
rect 519634 126511 519690 126520
rect 69018 125352 69074 125361
rect 69018 125287 69074 125296
rect 69032 124234 69060 125287
rect 69020 124228 69072 124234
rect 69020 124170 69072 124176
rect 519542 115560 519598 115569
rect 519542 115495 519598 115504
rect 69018 114472 69074 114481
rect 69018 114407 69074 114416
rect 69032 113218 69060 114407
rect 69020 113212 69072 113218
rect 69020 113154 69072 113160
rect 3698 110664 3754 110673
rect 3698 110599 3754 110608
rect 69018 103592 69074 103601
rect 3792 103556 3844 103562
rect 69018 103527 69020 103536
rect 3792 103498 3844 103504
rect 69072 103527 69074 103536
rect 69020 103498 69072 103504
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3700 92540 3752 92546
rect 3700 92482 3752 92488
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3608 81456 3660 81462
rect 3608 81398 3660 81404
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3516 70440 3568 70446
rect 3516 70382 3568 70388
rect 3424 59424 3476 59430
rect 3424 59366 3476 59372
rect 3436 6497 3464 59366
rect 3528 19417 3556 70382
rect 3620 32473 3648 81398
rect 3712 45529 3740 92482
rect 3804 58585 3832 103498
rect 69018 92712 69074 92721
rect 69018 92647 69074 92656
rect 69032 92546 69060 92647
rect 69020 92540 69072 92546
rect 69020 92482 69072 92488
rect 69018 81832 69074 81841
rect 69018 81767 69074 81776
rect 69032 81462 69060 81767
rect 69020 81456 69072 81462
rect 69020 81398 69072 81404
rect 519556 73166 519584 115495
rect 519648 86970 519676 126511
rect 519740 100706 519768 137663
rect 519832 113150 519860 148679
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 519820 113144 519872 113150
rect 519820 113086 519872 113092
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 519910 104408 519966 104417
rect 519910 104343 519966 104352
rect 519728 100700 519780 100706
rect 519728 100642 519780 100648
rect 519818 93256 519874 93265
rect 519818 93191 519874 93200
rect 519636 86964 519688 86970
rect 519636 86906 519688 86912
rect 519726 82240 519782 82249
rect 519726 82175 519782 82184
rect 519544 73160 519596 73166
rect 519544 73102 519596 73108
rect 519634 71088 519690 71097
rect 519634 71023 519690 71032
rect 69018 70816 69074 70825
rect 69018 70751 69074 70760
rect 69032 70446 69060 70751
rect 69020 70440 69072 70446
rect 69020 70382 69072 70388
rect 519542 60480 519598 60489
rect 519542 60415 519598 60424
rect 69018 60208 69074 60217
rect 69018 60143 69074 60152
rect 69032 59430 69060 60143
rect 72486 59922 72514 60044
rect 72436 59894 72514 59922
rect 69020 59424 69072 59430
rect 69020 59366 69072 59372
rect 3790 58576 3846 58585
rect 3790 58511 3846 58520
rect 72436 57934 72464 59894
rect 72886 59786 72914 60044
rect 72712 59758 72914 59786
rect 73786 59786 73814 60044
rect 74686 59786 74714 60044
rect 75586 59786 75614 60044
rect 76486 59786 76514 60044
rect 77386 59786 77414 60044
rect 73786 59758 73844 59786
rect 72424 57928 72476 57934
rect 72424 57870 72476 57876
rect 57244 57860 57296 57866
rect 57244 57802 57296 57808
rect 54484 57792 54536 57798
rect 54484 57734 54536 57740
rect 50344 57724 50396 57730
rect 50344 57666 50396 57672
rect 11704 57588 11756 57594
rect 11704 57530 11756 57536
rect 7564 57248 7616 57254
rect 7564 57190 7616 57196
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3606 32464 3662 32473
rect 3606 32399 3662 32408
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 6258
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 480 4108 3470
rect 5262 3360 5318 3369
rect 7576 3330 7604 57190
rect 7656 4956 7708 4962
rect 7656 4898 7708 4904
rect 5262 3295 5318 3304
rect 6460 3324 6512 3330
rect 5276 480 5304 3295
rect 6460 3266 6512 3272
rect 7564 3324 7616 3330
rect 7564 3266 7616 3272
rect 6472 480 6500 3266
rect 7668 480 7696 4898
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8772 480 8800 4762
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9968 480 9996 3538
rect 11150 3496 11206 3505
rect 11716 3466 11744 57530
rect 14464 57520 14516 57526
rect 14464 57462 14516 57468
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 11150 3431 11206 3440
rect 11704 3460 11756 3466
rect 11164 480 11192 3431
rect 11704 3402 11756 3408
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12360 480 12388 3062
rect 13556 480 13584 3606
rect 14476 3126 14504 57462
rect 18604 57452 18656 57458
rect 18604 57394 18656 57400
rect 15844 54528 15896 54534
rect 15844 54470 15896 54476
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14752 480 14780 3946
rect 15856 3602 15884 54470
rect 17868 13116 17920 13122
rect 17868 13058 17920 13064
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 17880 3534 17908 13058
rect 18616 4010 18644 57394
rect 29644 57384 29696 57390
rect 29644 57326 29696 57332
rect 22744 57316 22796 57322
rect 22744 57258 22796 57264
rect 22008 56160 22060 56166
rect 22008 56102 22060 56108
rect 22020 6914 22048 56102
rect 21836 6886 22048 6914
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18236 3800 18288 3806
rect 18236 3742 18288 3748
rect 19430 3768 19486 3777
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 480 15976 3334
rect 17052 480 17080 3470
rect 18248 480 18276 3742
rect 19430 3703 19486 3712
rect 19444 480 19472 3703
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 20640 480 20668 3567
rect 21836 480 21864 6886
rect 22756 3398 22784 57258
rect 25504 56024 25556 56030
rect 25504 55966 25556 55972
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 23032 480 23060 6122
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3538
rect 25516 3534 25544 55966
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 26528 480 26556 5034
rect 27724 480 27752 6190
rect 29656 3602 29684 57326
rect 41328 56364 41380 56370
rect 41328 56306 41380 56312
rect 37188 56296 37240 56302
rect 37188 56238 37240 56244
rect 34428 56228 34480 56234
rect 34428 56170 34480 56176
rect 32404 17264 32456 17270
rect 32404 17206 32456 17212
rect 31300 3868 31352 3874
rect 31300 3810 31352 3816
rect 29644 3596 29696 3602
rect 29644 3538 29696 3544
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 30116 480 30144 3062
rect 31312 480 31340 3810
rect 32416 3126 32444 17206
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32508 1850 32536 3538
rect 34440 3534 34468 56170
rect 35164 54596 35216 54602
rect 35164 54538 35216 54544
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 32416 1822 32536 1850
rect 32416 480 32444 1822
rect 33612 480 33640 3470
rect 34808 480 34836 4966
rect 35176 3670 35204 54538
rect 35164 3664 35216 3670
rect 35164 3606 35216 3612
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 36004 480 36032 3606
rect 37200 480 37228 56238
rect 39304 54664 39356 54670
rect 39304 54606 39356 54612
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 38396 480 38424 3878
rect 39316 3806 39344 54606
rect 39304 3800 39356 3806
rect 39304 3742 39356 3748
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39592 480 39620 3674
rect 41340 3398 41368 56306
rect 43444 56092 43496 56098
rect 43444 56034 43496 56040
rect 42984 7608 43036 7614
rect 42984 7550 43036 7556
rect 42996 3398 43024 7550
rect 43456 3874 43484 56034
rect 47584 54732 47636 54738
rect 47584 54674 47636 54680
rect 44272 5160 44324 5166
rect 44272 5102 44324 5108
rect 43444 3868 43496 3874
rect 43444 3810 43496 3816
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3334
rect 43088 480 43116 3742
rect 44284 480 44312 5102
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45480 480 45508 4014
rect 47596 3942 47624 54674
rect 47860 8968 47912 8974
rect 47860 8910 47912 8916
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 46664 3868 46716 3874
rect 46664 3810 46716 3816
rect 46676 480 46704 3810
rect 47872 480 47900 8910
rect 50356 5030 50384 57666
rect 53104 57656 53156 57662
rect 53104 57598 53156 57604
rect 51724 25560 51776 25566
rect 51724 25502 51776 25508
rect 50344 5024 50396 5030
rect 50344 4966 50396 4972
rect 48964 4208 49016 4214
rect 48964 4150 49016 4156
rect 48976 480 49004 4150
rect 51736 4078 51764 25502
rect 52368 15904 52420 15910
rect 52368 15846 52420 15852
rect 51724 4072 51776 4078
rect 51724 4014 51776 4020
rect 50160 4004 50212 4010
rect 50160 3946 50212 3952
rect 50172 480 50200 3946
rect 52380 3398 52408 15846
rect 52552 8288 52604 8294
rect 52552 8230 52604 8236
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 51368 480 51396 3334
rect 52564 480 52592 8230
rect 53116 4214 53144 57598
rect 54496 8294 54524 57734
rect 54944 14476 54996 14482
rect 54944 14418 54996 14424
rect 54484 8288 54536 8294
rect 54484 8230 54536 8236
rect 53104 4208 53156 4214
rect 53104 4150 53156 4156
rect 53748 4140 53800 4146
rect 53748 4082 53800 4088
rect 53760 480 53788 4082
rect 54956 480 54984 14418
rect 57256 5098 57284 57802
rect 71044 57588 71096 57594
rect 71044 57530 71096 57536
rect 68284 57180 68336 57186
rect 68284 57122 68336 57128
rect 65616 56976 65668 56982
rect 65616 56918 65668 56924
rect 62028 56432 62080 56438
rect 62028 56374 62080 56380
rect 58624 55888 58676 55894
rect 58624 55830 58676 55836
rect 57336 11824 57388 11830
rect 57336 11766 57388 11772
rect 57244 5092 57296 5098
rect 57244 5034 57296 5040
rect 56048 5024 56100 5030
rect 56048 4966 56100 4972
rect 56060 480 56088 4966
rect 57348 4146 57376 11766
rect 57336 4140 57388 4146
rect 57336 4082 57388 4088
rect 58636 4010 58664 55830
rect 61936 29640 61988 29646
rect 61936 29582 61988 29588
rect 59268 19984 59320 19990
rect 59268 19926 59320 19932
rect 58624 4004 58676 4010
rect 58624 3946 58676 3952
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 57256 480 57284 3878
rect 59280 3398 59308 19926
rect 59636 5228 59688 5234
rect 59636 5170 59688 5176
rect 58440 3392 58492 3398
rect 58440 3334 58492 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 58452 480 58480 3334
rect 59648 480 59676 5170
rect 61948 3398 61976 29582
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 61936 3392 61988 3398
rect 61936 3334 61988 3340
rect 60844 480 60872 3334
rect 62040 480 62068 56374
rect 65524 55956 65576 55962
rect 65524 55898 65576 55904
rect 65536 6914 65564 55898
rect 65628 14482 65656 56918
rect 68296 15910 68324 57122
rect 69664 57112 69716 57118
rect 69664 57054 69716 57060
rect 68376 18624 68428 18630
rect 68376 18566 68428 18572
rect 68284 15904 68336 15910
rect 68284 15846 68336 15852
rect 65616 14476 65668 14482
rect 65616 14418 65668 14424
rect 66168 10328 66220 10334
rect 66168 10270 66220 10276
rect 65444 6886 65564 6914
rect 63224 6384 63276 6390
rect 63224 6326 63276 6332
rect 63236 480 63264 6326
rect 65444 4146 65472 6886
rect 64328 4140 64380 4146
rect 64328 4082 64380 4088
rect 65432 4140 65484 4146
rect 65432 4082 65484 4088
rect 64340 480 64368 4082
rect 66180 3398 66208 10270
rect 66720 5092 66772 5098
rect 66720 5034 66772 5040
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 66168 3392 66220 3398
rect 66168 3334 66220 3340
rect 65536 480 65564 3334
rect 66732 480 66760 5034
rect 68388 3942 68416 18566
rect 69676 9042 69704 57054
rect 69664 9036 69716 9042
rect 69664 8978 69716 8984
rect 69112 8968 69164 8974
rect 69112 8910 69164 8916
rect 68376 3936 68428 3942
rect 68376 3878 68428 3884
rect 67916 3052 67968 3058
rect 67916 2994 67968 3000
rect 67928 480 67956 2994
rect 69124 480 69152 8910
rect 70308 7676 70360 7682
rect 70308 7618 70360 7624
rect 70320 480 70348 7618
rect 71056 6322 71084 57530
rect 71780 57044 71832 57050
rect 71780 56986 71832 56992
rect 71792 56370 71820 56986
rect 71780 56364 71832 56370
rect 71780 56306 71832 56312
rect 72712 45554 72740 59758
rect 73816 57594 73844 59758
rect 74644 59758 74714 59786
rect 75564 59758 75614 59786
rect 75932 59758 76514 59786
rect 77312 59758 77414 59786
rect 78306 59786 78334 60044
rect 79206 59786 79234 60044
rect 80106 59786 80134 60044
rect 81006 59786 81034 60044
rect 78306 59758 78352 59786
rect 73804 57588 73856 57594
rect 73804 57530 73856 57536
rect 71884 45526 72740 45554
rect 71044 6316 71096 6322
rect 71044 6258 71096 6264
rect 71228 6316 71280 6322
rect 71228 6258 71280 6264
rect 71240 3058 71268 6258
rect 71884 4894 71912 45526
rect 72608 5296 72660 5302
rect 72608 5238 72660 5244
rect 71872 4888 71924 4894
rect 71872 4830 71924 4836
rect 71504 4140 71556 4146
rect 71504 4082 71556 4088
rect 71228 3052 71280 3058
rect 71228 2994 71280 3000
rect 71516 480 71544 4082
rect 72620 480 72648 5238
rect 74644 4962 74672 59758
rect 75564 57526 75592 59758
rect 75552 57520 75604 57526
rect 75552 57462 75604 57468
rect 75828 57520 75880 57526
rect 75828 57462 75880 57468
rect 74632 4956 74684 4962
rect 74632 4898 74684 4904
rect 73804 4888 73856 4894
rect 73804 4830 73856 4836
rect 73816 480 73844 4830
rect 75840 3398 75868 57462
rect 75932 13122 75960 59758
rect 77312 56658 77340 59758
rect 78324 57866 78352 59758
rect 78692 59758 79234 59786
rect 80072 59758 80134 59786
rect 80992 59758 81034 59786
rect 81906 59786 81934 60044
rect 82806 59786 82834 60044
rect 83706 59786 83734 60044
rect 84626 59786 84654 60044
rect 85526 59786 85554 60044
rect 86426 59786 86454 60044
rect 81906 59758 81940 59786
rect 82806 59758 82860 59786
rect 78312 57860 78364 57866
rect 78312 57802 78364 57808
rect 77220 56630 77340 56658
rect 77220 56166 77248 56630
rect 77208 56160 77260 56166
rect 77208 56102 77260 56108
rect 78692 17270 78720 59758
rect 79324 57588 79376 57594
rect 79324 57530 79376 57536
rect 78680 17264 78732 17270
rect 78680 17206 78732 17212
rect 75920 13116 75972 13122
rect 75920 13058 75972 13064
rect 76564 13116 76616 13122
rect 76564 13058 76616 13064
rect 76196 5364 76248 5370
rect 76196 5306 76248 5312
rect 75000 3392 75052 3398
rect 75000 3334 75052 3340
rect 75828 3392 75880 3398
rect 75828 3334 75880 3340
rect 75012 480 75040 3334
rect 76208 480 76236 5306
rect 76576 4146 76604 13058
rect 79336 5234 79364 57530
rect 80072 56658 80100 59758
rect 79980 56630 80100 56658
rect 79980 56234 80008 56630
rect 80992 56302 81020 59758
rect 81912 57050 81940 59758
rect 81900 57044 81952 57050
rect 81900 56986 81952 56992
rect 80980 56296 81032 56302
rect 80980 56238 81032 56244
rect 79968 56228 80020 56234
rect 79968 56170 80020 56176
rect 81348 24132 81400 24138
rect 81348 24074 81400 24080
rect 79324 5228 79376 5234
rect 79324 5170 79376 5176
rect 79692 5228 79744 5234
rect 79692 5170 79744 5176
rect 77392 4956 77444 4962
rect 77392 4898 77444 4904
rect 76564 4140 76616 4146
rect 76564 4082 76616 4088
rect 77404 480 77432 4898
rect 78588 3936 78640 3942
rect 78588 3878 78640 3884
rect 78600 480 78628 3878
rect 79704 480 79732 5170
rect 81360 3398 81388 24074
rect 82832 5166 82860 59758
rect 83660 59758 83734 59786
rect 84580 59758 84654 59786
rect 85500 59758 85554 59786
rect 85592 59758 86454 59786
rect 86960 59832 87012 59838
rect 86960 59774 87012 59780
rect 87326 59786 87354 60044
rect 88226 59838 88254 60044
rect 88214 59832 88266 59838
rect 83660 57118 83688 59758
rect 84580 57186 84608 59758
rect 85500 57934 85528 59758
rect 85488 57928 85540 57934
rect 85488 57870 85540 57876
rect 84568 57180 84620 57186
rect 84568 57122 84620 57128
rect 83648 57112 83700 57118
rect 83648 57054 83700 57060
rect 85592 19990 85620 59758
rect 86224 56840 86276 56846
rect 86224 56782 86276 56788
rect 85580 19984 85632 19990
rect 85580 19926 85632 19932
rect 83280 5432 83332 5438
rect 83280 5374 83332 5380
rect 82820 5160 82872 5166
rect 82820 5102 82872 5108
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3946
rect 83292 480 83320 5374
rect 86236 5302 86264 56782
rect 86972 10334 87000 59774
rect 87326 59758 87368 59786
rect 89126 59786 89154 60044
rect 88214 59774 88266 59780
rect 87340 56438 87368 59758
rect 88352 59758 89154 59786
rect 89812 59832 89864 59838
rect 90046 59786 90074 60044
rect 90946 59838 90974 60044
rect 89812 59774 89864 59780
rect 87604 57928 87656 57934
rect 87604 57870 87656 57876
rect 87328 56432 87380 56438
rect 87328 56374 87380 56380
rect 86960 10328 87012 10334
rect 86960 10270 87012 10276
rect 87616 5438 87644 57870
rect 88352 8974 88380 59758
rect 88984 57860 89036 57866
rect 88984 57802 89036 57808
rect 88340 8968 88392 8974
rect 88340 8910 88392 8916
rect 87972 6452 88024 6458
rect 87972 6394 88024 6400
rect 87604 5432 87656 5438
rect 87604 5374 87656 5380
rect 86224 5296 86276 5302
rect 86224 5238 86276 5244
rect 84476 5160 84528 5166
rect 84476 5102 84528 5108
rect 84488 480 84516 5102
rect 86868 4208 86920 4214
rect 86868 4150 86920 4156
rect 85672 4072 85724 4078
rect 85672 4014 85724 4020
rect 85684 480 85712 4014
rect 86880 480 86908 4150
rect 87984 480 88012 6394
rect 88996 5234 89024 57802
rect 89824 5370 89852 59774
rect 90008 59758 90074 59786
rect 90934 59832 90986 59838
rect 90934 59774 90986 59780
rect 91846 59786 91874 60044
rect 92746 59922 92774 60044
rect 92492 59894 92774 59922
rect 91846 59758 91876 59786
rect 90008 56846 90036 59758
rect 91848 57866 91876 59758
rect 92492 57934 92520 59894
rect 93646 59786 93674 60044
rect 94546 59786 94574 60044
rect 95446 59786 95474 60044
rect 92584 59758 93674 59786
rect 93872 59758 94574 59786
rect 95252 59758 95474 59786
rect 96366 59786 96394 60044
rect 97266 59786 97294 60044
rect 98166 59786 98194 60044
rect 99066 59786 99094 60044
rect 99966 59786 99994 60044
rect 100866 59786 100894 60044
rect 96366 59758 96568 59786
rect 97266 59758 97304 59786
rect 98166 59758 98224 59786
rect 99066 59758 99328 59786
rect 92480 57928 92532 57934
rect 92480 57870 92532 57876
rect 91836 57860 91888 57866
rect 91836 57802 91888 57808
rect 89996 56840 90048 56846
rect 89996 56782 90048 56788
rect 89812 5364 89864 5370
rect 89812 5306 89864 5312
rect 88984 5228 89036 5234
rect 88984 5170 89036 5176
rect 91560 5228 91612 5234
rect 91560 5170 91612 5176
rect 90364 4548 90416 4554
rect 90364 4490 90416 4496
rect 89168 4140 89220 4146
rect 89168 4082 89220 4088
rect 89180 480 89208 4082
rect 90376 480 90404 4490
rect 91572 480 91600 5170
rect 92584 4214 92612 59758
rect 93872 4554 93900 59758
rect 95252 57610 95280 59758
rect 95160 57582 95280 57610
rect 96540 57610 96568 59758
rect 97276 57866 97304 59758
rect 98196 57866 98224 59758
rect 97264 57860 97316 57866
rect 97264 57802 97316 57808
rect 97908 57860 97960 57866
rect 97908 57802 97960 57808
rect 98184 57860 98236 57866
rect 98184 57802 98236 57808
rect 99196 57860 99248 57866
rect 99196 57802 99248 57808
rect 96540 57582 96660 57610
rect 95056 6520 95108 6526
rect 95056 6462 95108 6468
rect 93860 4548 93912 4554
rect 93860 4490 93912 4496
rect 92572 4208 92624 4214
rect 92572 4150 92624 4156
rect 92756 3392 92808 3398
rect 92756 3334 92808 3340
rect 92768 480 92796 3334
rect 93952 3324 94004 3330
rect 93952 3266 94004 3272
rect 93964 480 93992 3266
rect 95068 3210 95096 6462
rect 95160 3330 95188 57582
rect 96632 16574 96660 57582
rect 96632 16546 97488 16574
rect 95148 3324 95200 3330
rect 95148 3266 95200 3272
rect 96252 3256 96304 3262
rect 95068 3182 95188 3210
rect 96252 3198 96304 3204
rect 95160 480 95188 3182
rect 96264 480 96292 3198
rect 97460 480 97488 16546
rect 97920 4214 97948 57802
rect 98644 6588 98696 6594
rect 98644 6530 98696 6536
rect 97908 4208 97960 4214
rect 97908 4150 97960 4156
rect 98656 480 98684 6530
rect 99208 4622 99236 57802
rect 99300 4758 99328 59758
rect 99944 59758 99994 59786
rect 100864 59758 100894 59786
rect 101766 59786 101794 60044
rect 102686 59786 102714 60044
rect 103586 59786 103614 60044
rect 104486 59786 104514 60044
rect 105386 59786 105414 60044
rect 101766 59758 101996 59786
rect 102686 59758 102732 59786
rect 99944 57866 99972 59758
rect 100668 57928 100720 57934
rect 100668 57870 100720 57876
rect 99932 57860 99984 57866
rect 99932 57802 99984 57808
rect 100576 57860 100628 57866
rect 100576 57802 100628 57808
rect 100588 5506 100616 57802
rect 100576 5500 100628 5506
rect 100576 5442 100628 5448
rect 99288 4752 99340 4758
rect 99288 4694 99340 4700
rect 99196 4616 99248 4622
rect 99196 4558 99248 4564
rect 100680 3330 100708 57870
rect 100864 57866 100892 59758
rect 100852 57860 100904 57866
rect 100852 57802 100904 57808
rect 101968 5302 101996 59758
rect 102048 57860 102100 57866
rect 102048 57802 102100 57808
rect 102060 5438 102088 57802
rect 102704 56642 102732 59758
rect 103532 59758 103614 59786
rect 103716 59758 104514 59786
rect 104912 59758 105414 59786
rect 106286 59786 106314 60044
rect 107186 59786 107214 60044
rect 108106 59786 108134 60044
rect 106286 59758 106412 59786
rect 102692 56636 102744 56642
rect 102692 56578 102744 56584
rect 103532 56030 103560 59758
rect 103520 56024 103572 56030
rect 103520 55966 103572 55972
rect 102232 6656 102284 6662
rect 102232 6598 102284 6604
rect 102048 5432 102100 5438
rect 102048 5374 102100 5380
rect 101956 5296 102008 5302
rect 101956 5238 102008 5244
rect 101036 4208 101088 4214
rect 101036 4150 101088 4156
rect 99840 3324 99892 3330
rect 99840 3266 99892 3272
rect 100668 3324 100720 3330
rect 100668 3266 100720 3272
rect 99852 480 99880 3266
rect 101048 480 101076 4150
rect 102244 480 102272 6598
rect 103716 4826 103744 59758
rect 104912 54602 104940 59758
rect 106280 57724 106332 57730
rect 106280 57666 106332 57672
rect 105544 56636 105596 56642
rect 105544 56578 105596 56584
rect 104900 54596 104952 54602
rect 104900 54538 104952 54544
rect 105556 5370 105584 56578
rect 105728 8968 105780 8974
rect 105728 8910 105780 8916
rect 105544 5364 105596 5370
rect 105544 5306 105596 5312
rect 103704 4820 103756 4826
rect 103704 4762 103756 4768
rect 104532 4616 104584 4622
rect 104532 4558 104584 4564
rect 103336 3256 103388 3262
rect 103336 3198 103388 3204
rect 103348 480 103376 3198
rect 104544 480 104572 4558
rect 105740 480 105768 8910
rect 106292 6186 106320 57666
rect 106384 54670 106412 59758
rect 107120 59758 107214 59786
rect 107672 59758 108134 59786
rect 109006 59786 109034 60044
rect 109906 59786 109934 60044
rect 109006 59758 109080 59786
rect 107120 57730 107148 59758
rect 107108 57724 107160 57730
rect 107108 57666 107160 57672
rect 106372 54664 106424 54670
rect 106372 54606 106424 54612
rect 107672 6254 107700 59758
rect 109052 56098 109080 59758
rect 109880 59758 109934 59786
rect 110420 59832 110472 59838
rect 110806 59786 110834 60044
rect 111706 59838 111734 60044
rect 110420 59774 110472 59780
rect 109880 57934 109908 59758
rect 109868 57928 109920 57934
rect 109868 57870 109920 57876
rect 109040 56092 109092 56098
rect 109040 56034 109092 56040
rect 110432 7614 110460 59774
rect 110524 59758 110834 59786
rect 111694 59832 111746 59838
rect 112606 59786 112634 60044
rect 113506 59786 113534 60044
rect 114426 59786 114454 60044
rect 115326 59786 115354 60044
rect 116226 59922 116254 60044
rect 111694 59774 111746 59780
rect 111812 59758 112634 59786
rect 113468 59758 113534 59786
rect 114388 59758 114454 59786
rect 114664 59758 115354 59786
rect 115952 59894 116254 59922
rect 110524 54738 110552 59758
rect 110512 54732 110564 54738
rect 110512 54674 110564 54680
rect 111812 25566 111840 59758
rect 113468 57662 113496 59758
rect 114388 57798 114416 59758
rect 114376 57792 114428 57798
rect 114376 57734 114428 57740
rect 113456 57656 113508 57662
rect 113456 57598 113508 57604
rect 111800 25560 111852 25566
rect 111800 25502 111852 25508
rect 113088 25560 113140 25566
rect 113088 25502 113140 25508
rect 110420 7608 110472 7614
rect 110420 7550 110472 7556
rect 113100 6914 113128 25502
rect 112824 6886 113128 6914
rect 107660 6248 107712 6254
rect 107660 6190 107712 6196
rect 106280 6180 106332 6186
rect 106280 6122 106332 6128
rect 111616 5500 111668 5506
rect 111616 5442 111668 5448
rect 109316 4820 109368 4826
rect 109316 4762 109368 4768
rect 108120 4752 108172 4758
rect 108120 4694 108172 4700
rect 106924 3188 106976 3194
rect 106924 3130 106976 3136
rect 106936 480 106964 3130
rect 108132 480 108160 4694
rect 109328 480 109356 4762
rect 110512 3120 110564 3126
rect 110512 3062 110564 3068
rect 110524 480 110552 3062
rect 111628 480 111656 5442
rect 112824 480 112852 6886
rect 114664 5030 114692 59758
rect 115204 57724 115256 57730
rect 115204 57666 115256 57672
rect 115112 5432 115164 5438
rect 115112 5374 115164 5380
rect 114652 5024 114704 5030
rect 114652 4966 114704 4972
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114020 480 114048 2994
rect 115124 2802 115152 5374
rect 115216 4962 115244 57666
rect 115952 57594 115980 59894
rect 117126 59786 117154 60044
rect 118026 59786 118054 60044
rect 118926 59786 118954 60044
rect 119826 59786 119854 60044
rect 120746 59786 120774 60044
rect 121646 59786 121674 60044
rect 122546 59786 122574 60044
rect 123446 59786 123474 60044
rect 124346 59786 124374 60044
rect 125246 59786 125274 60044
rect 126166 59786 126194 60044
rect 116044 59758 117154 59786
rect 117976 59758 118054 59786
rect 118712 59758 118954 59786
rect 119080 59758 119854 59786
rect 120736 59758 120774 59786
rect 121472 59758 121674 59786
rect 121748 59758 122574 59786
rect 122852 59758 123474 59786
rect 124324 59758 124374 59786
rect 124416 59758 125274 59786
rect 125612 59758 126194 59786
rect 127066 59786 127094 60044
rect 127966 59786 127994 60044
rect 128866 59786 128894 60044
rect 127066 59758 127112 59786
rect 115940 57588 115992 57594
rect 115940 57530 115992 57536
rect 116044 6390 116072 59758
rect 117976 57662 118004 59758
rect 116584 57656 116636 57662
rect 116584 57598 116636 57604
rect 117964 57656 118016 57662
rect 117964 57598 118016 57604
rect 116032 6384 116084 6390
rect 116032 6326 116084 6332
rect 116400 6248 116452 6254
rect 116400 6190 116452 6196
rect 115204 4956 115256 4962
rect 115204 4898 115256 4904
rect 115124 2774 115244 2802
rect 115216 480 115244 2774
rect 116412 480 116440 6190
rect 116596 5098 116624 57598
rect 118712 7682 118740 59758
rect 119080 45554 119108 59758
rect 120736 57730 120764 59758
rect 120724 57724 120776 57730
rect 120724 57666 120776 57672
rect 118896 45526 119108 45554
rect 118700 7676 118752 7682
rect 118700 7618 118752 7624
rect 118792 5296 118844 5302
rect 118792 5238 118844 5244
rect 116584 5092 116636 5098
rect 116584 5034 116636 5040
rect 117596 2984 117648 2990
rect 117596 2926 117648 2932
rect 117608 480 117636 2926
rect 118804 480 118832 5238
rect 118896 4894 118924 45526
rect 121472 24138 121500 59758
rect 121748 45554 121776 59758
rect 121656 45526 121776 45554
rect 121460 24132 121512 24138
rect 121460 24074 121512 24080
rect 119896 7608 119948 7614
rect 119896 7550 119948 7556
rect 118884 4888 118936 4894
rect 118884 4830 118936 4836
rect 119908 480 119936 7550
rect 121656 5166 121684 45526
rect 122852 6458 122880 59758
rect 124324 57662 124352 59758
rect 123484 57656 123536 57662
rect 123484 57598 123536 57604
rect 124312 57656 124364 57662
rect 124312 57598 124364 57604
rect 122840 6452 122892 6458
rect 122840 6394 122892 6400
rect 122288 5364 122340 5370
rect 122288 5306 122340 5312
rect 121644 5160 121696 5166
rect 121644 5102 121696 5108
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 5306
rect 123496 5234 123524 57598
rect 124416 45554 124444 59758
rect 124864 57588 124916 57594
rect 124864 57530 124916 57536
rect 124324 45526 124444 45554
rect 124324 6526 124352 45526
rect 124876 8974 124904 57530
rect 124864 8968 124916 8974
rect 124864 8910 124916 8916
rect 125612 6594 125640 59758
rect 127084 57662 127112 59758
rect 127912 59758 127994 59786
rect 128372 59758 128894 59786
rect 129766 59786 129794 60044
rect 130666 59786 130694 60044
rect 131566 59786 131594 60044
rect 132486 59786 132514 60044
rect 133386 59786 133414 60044
rect 129766 59758 129872 59786
rect 130666 59758 130700 59786
rect 131566 59758 131620 59786
rect 132486 59758 132540 59786
rect 126244 57656 126296 57662
rect 126244 57598 126296 57604
rect 127072 57656 127124 57662
rect 127072 57598 127124 57604
rect 126256 6662 126284 57598
rect 127912 57594 127940 59758
rect 127900 57588 127952 57594
rect 127900 57530 127952 57536
rect 128176 10328 128228 10334
rect 128176 10270 128228 10276
rect 126980 7064 127032 7070
rect 126980 7006 127032 7012
rect 126244 6656 126296 6662
rect 126244 6598 126296 6604
rect 125600 6588 125652 6594
rect 125600 6530 125652 6536
rect 124312 6520 124364 6526
rect 124312 6462 124364 6468
rect 125876 6180 125928 6186
rect 125876 6122 125928 6128
rect 123484 5228 123536 5234
rect 123484 5170 123536 5176
rect 123484 4888 123536 4894
rect 123484 4830 123536 4836
rect 123496 480 123524 4830
rect 124680 2848 124732 2854
rect 124680 2790 124732 2796
rect 124692 480 124720 2790
rect 125888 480 125916 6122
rect 126992 480 127020 7006
rect 128188 480 128216 10270
rect 128372 4826 128400 59758
rect 129740 57656 129792 57662
rect 129740 57598 129792 57604
rect 129004 57588 129056 57594
rect 129004 57530 129056 57536
rect 129016 7614 129044 57530
rect 129004 7608 129056 7614
rect 129004 7550 129056 7556
rect 129752 6254 129780 57598
rect 129844 25566 129872 59758
rect 130672 57662 130700 59758
rect 130660 57656 130712 57662
rect 130660 57598 130712 57604
rect 131592 57594 131620 59758
rect 131580 57588 131632 57594
rect 131580 57530 131632 57536
rect 129832 25560 129884 25566
rect 129832 25502 129884 25508
rect 131764 10396 131816 10402
rect 131764 10338 131816 10344
rect 130568 8968 130620 8974
rect 130568 8910 130620 8916
rect 129740 6248 129792 6254
rect 129740 6190 129792 6196
rect 128360 4820 128412 4826
rect 128360 4762 128412 4768
rect 129372 4820 129424 4826
rect 129372 4762 129424 4768
rect 129384 480 129412 4762
rect 130580 480 130608 8910
rect 131776 480 131804 10338
rect 132512 4894 132540 59758
rect 132604 59758 133414 59786
rect 133972 59832 134024 59838
rect 134286 59786 134314 60044
rect 135186 59838 135214 60044
rect 133972 59774 134024 59780
rect 132604 54534 132632 59758
rect 132592 54528 132644 54534
rect 132592 54470 132644 54476
rect 132500 4888 132552 4894
rect 132500 4830 132552 4836
rect 132960 4888 133012 4894
rect 132960 4830 133012 4836
rect 132972 480 133000 4830
rect 133984 3777 134012 59774
rect 134260 59758 134314 59786
rect 135174 59832 135226 59838
rect 136086 59786 136114 60044
rect 135174 59774 135226 59780
rect 135456 59758 136114 59786
rect 136640 59832 136692 59838
rect 136986 59786 137014 60044
rect 137886 59838 137914 60044
rect 136640 59774 136692 59780
rect 134260 57458 134288 59758
rect 134248 57452 134300 57458
rect 134248 57394 134300 57400
rect 134156 9036 134208 9042
rect 134156 8978 134208 8984
rect 133970 3768 134026 3777
rect 133970 3703 134026 3712
rect 134168 480 134196 8978
rect 135260 3528 135312 3534
rect 135260 3470 135312 3476
rect 135272 480 135300 3470
rect 135456 3466 135484 59758
rect 136456 11756 136508 11762
rect 136456 11698 136508 11704
rect 136468 3534 136496 11698
rect 136548 4956 136600 4962
rect 136548 4898 136600 4904
rect 136456 3528 136508 3534
rect 136456 3470 136508 3476
rect 135444 3460 135496 3466
rect 135444 3402 135496 3408
rect 136560 2530 136588 4898
rect 136652 3602 136680 59774
rect 136836 59758 137014 59786
rect 137874 59832 137926 59838
rect 138806 59786 138834 60044
rect 137874 59774 137926 59780
rect 138032 59758 138834 59786
rect 139400 59832 139452 59838
rect 139706 59786 139734 60044
rect 140606 59838 140634 60044
rect 139400 59774 139452 59780
rect 136836 3738 136864 59758
rect 137652 14748 137704 14754
rect 137652 14690 137704 14696
rect 136824 3732 136876 3738
rect 136824 3674 136876 3680
rect 136640 3596 136692 3602
rect 136640 3538 136692 3544
rect 136468 2502 136588 2530
rect 136468 480 136496 2502
rect 137664 480 137692 14690
rect 138032 3670 138060 59758
rect 139308 15904 139360 15910
rect 139308 15846 139360 15852
rect 138020 3664 138072 3670
rect 138020 3606 138072 3612
rect 139320 3534 139348 15846
rect 139412 3806 139440 59774
rect 139504 59758 139734 59786
rect 140594 59832 140646 59838
rect 141506 59786 141534 60044
rect 140594 59774 140646 59780
rect 140792 59758 141534 59786
rect 142160 59832 142212 59838
rect 142406 59786 142434 60044
rect 143306 59838 143334 60044
rect 142160 59774 142212 59780
rect 139400 3800 139452 3806
rect 139400 3742 139452 3748
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 138860 480 138888 3470
rect 139504 3466 139532 59758
rect 140044 5092 140096 5098
rect 140044 5034 140096 5040
rect 139492 3460 139544 3466
rect 139492 3402 139544 3408
rect 140056 480 140084 5034
rect 140792 3874 140820 59758
rect 142068 36576 142120 36582
rect 142068 36518 142120 36524
rect 140780 3868 140832 3874
rect 140780 3810 140832 3816
rect 142080 3534 142108 36518
rect 142172 11830 142200 59774
rect 142356 59758 142434 59786
rect 143294 59832 143346 59838
rect 144226 59786 144254 60044
rect 145126 59786 145154 60044
rect 143294 59774 143346 59780
rect 143552 59758 144254 59786
rect 145116 59758 145154 59786
rect 146026 59786 146054 60044
rect 146926 59786 146954 60044
rect 147826 59786 147854 60044
rect 148726 59786 148754 60044
rect 149626 59786 149654 60044
rect 146026 59758 146064 59786
rect 142356 55894 142384 59758
rect 142344 55888 142396 55894
rect 142344 55830 142396 55836
rect 143552 18630 143580 59758
rect 145116 57662 145144 59758
rect 144184 57656 144236 57662
rect 144184 57598 144236 57604
rect 145104 57656 145156 57662
rect 145104 57598 145156 57604
rect 144196 29646 144224 57598
rect 146036 55962 146064 59758
rect 146312 59758 146954 59786
rect 147784 59758 147854 59786
rect 148704 59758 148754 59786
rect 149072 59758 149654 59786
rect 150440 59832 150492 59838
rect 150546 59786 150574 60044
rect 151446 59838 151474 60044
rect 150440 59774 150492 59780
rect 146024 55956 146076 55962
rect 146024 55898 146076 55904
rect 144184 29640 144236 29646
rect 144184 29582 144236 29588
rect 144828 28280 144880 28286
rect 144828 28222 144880 28228
rect 143540 18624 143592 18630
rect 143540 18566 143592 18572
rect 143448 17264 143500 17270
rect 143448 17206 143500 17212
rect 142160 11824 142212 11830
rect 142160 11766 142212 11772
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 141252 480 141280 3470
rect 143460 3466 143488 17206
rect 144736 14816 144788 14822
rect 144736 14758 144788 14764
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 142436 3460 142488 3466
rect 142436 3402 142488 3408
rect 143448 3460 143500 3466
rect 143448 3402 143500 3408
rect 142448 480 142476 3402
rect 143552 480 143580 3470
rect 144748 480 144776 14758
rect 144840 3534 144868 28222
rect 146312 6322 146340 59758
rect 147784 13122 147812 59758
rect 148704 57526 148732 59758
rect 148968 57588 149020 57594
rect 148968 57530 149020 57536
rect 148692 57520 148744 57526
rect 148692 57462 148744 57468
rect 147772 13116 147824 13122
rect 147772 13058 147824 13064
rect 146300 6316 146352 6322
rect 146300 6258 146352 6264
rect 147128 5024 147180 5030
rect 147128 4966 147180 4972
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 145932 3460 145984 3466
rect 145932 3402 145984 3408
rect 145944 480 145972 3402
rect 147140 480 147168 4966
rect 148980 3534 149008 57530
rect 149072 3942 149100 59758
rect 150452 4078 150480 59774
rect 150544 59758 150574 59786
rect 151434 59832 151486 59838
rect 152346 59786 152374 60044
rect 151434 59774 151486 59780
rect 151832 59758 152374 59786
rect 153246 59786 153274 60044
rect 154146 59786 154174 60044
rect 153246 59758 153332 59786
rect 150440 4072 150492 4078
rect 150440 4014 150492 4020
rect 150544 4010 150572 59758
rect 151832 4010 151860 59758
rect 153200 57656 153252 57662
rect 153200 57598 153252 57604
rect 153108 31068 153160 31074
rect 153108 31010 153160 31016
rect 150532 4004 150584 4010
rect 150532 3946 150584 3952
rect 151820 4004 151872 4010
rect 151820 3946 151872 3952
rect 149060 3936 149112 3942
rect 149060 3878 149112 3884
rect 150624 3800 150676 3806
rect 150624 3742 150676 3748
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 150636 480 150664 3742
rect 153120 3602 153148 31010
rect 151820 3596 151872 3602
rect 151820 3538 151872 3544
rect 153108 3596 153160 3602
rect 153108 3538 153160 3544
rect 151832 480 151860 3538
rect 153016 3392 153068 3398
rect 153016 3334 153068 3340
rect 153028 480 153056 3334
rect 153212 3262 153240 57598
rect 153304 3330 153332 59758
rect 154132 59758 154174 59786
rect 155046 59786 155074 60044
rect 155946 59786 155974 60044
rect 156866 59786 156894 60044
rect 155046 59758 155080 59786
rect 155946 59758 156000 59786
rect 154132 57662 154160 59758
rect 155052 57866 155080 59758
rect 155040 57860 155092 57866
rect 155040 57802 155092 57808
rect 155868 57724 155920 57730
rect 155868 57666 155920 57672
rect 154120 57656 154172 57662
rect 154120 57598 154172 57604
rect 154212 3868 154264 3874
rect 154212 3810 154264 3816
rect 153292 3324 153344 3330
rect 153292 3266 153344 3272
rect 153200 3256 153252 3262
rect 153200 3198 153252 3204
rect 154224 480 154252 3810
rect 155880 3602 155908 57666
rect 155408 3596 155460 3602
rect 155408 3538 155460 3544
rect 155868 3596 155920 3602
rect 155868 3538 155920 3544
rect 155420 480 155448 3538
rect 155972 3194 156000 59758
rect 156064 59758 156894 59786
rect 157340 59832 157392 59838
rect 157766 59786 157794 60044
rect 158666 59838 158694 60044
rect 157340 59774 157392 59780
rect 155960 3188 156012 3194
rect 155960 3130 156012 3136
rect 156064 3126 156092 59758
rect 156604 3664 156656 3670
rect 156604 3606 156656 3612
rect 156052 3120 156104 3126
rect 156052 3062 156104 3068
rect 156616 480 156644 3606
rect 157352 2990 157380 59774
rect 157444 59758 157794 59786
rect 158654 59832 158706 59838
rect 159566 59786 159594 60044
rect 158654 59774 158706 59780
rect 158824 59758 159594 59786
rect 160192 59832 160244 59838
rect 160466 59786 160494 60044
rect 161366 59838 161394 60044
rect 160192 59774 160244 59780
rect 157444 3058 157472 59758
rect 157800 3936 157852 3942
rect 157800 3878 157852 3884
rect 157432 3052 157484 3058
rect 157432 2994 157484 3000
rect 157340 2984 157392 2990
rect 157340 2926 157392 2932
rect 157812 480 157840 3878
rect 158824 2922 158852 59758
rect 160008 32428 160060 32434
rect 160008 32370 160060 32376
rect 160020 3602 160048 32370
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 158904 3596 158956 3602
rect 158904 3538 158956 3544
rect 160008 3596 160060 3602
rect 160008 3538 160060 3544
rect 158812 2916 158864 2922
rect 158812 2858 158864 2864
rect 158916 480 158944 3538
rect 160112 480 160140 3674
rect 160204 2854 160232 59774
rect 160388 59758 160494 59786
rect 161354 59832 161406 59838
rect 162286 59786 162314 60044
rect 161354 59774 161406 59780
rect 161584 59758 162314 59786
rect 162952 59832 163004 59838
rect 163186 59786 163214 60044
rect 164086 59838 164114 60044
rect 162952 59774 163004 59780
rect 160388 4010 160416 59758
rect 161388 57452 161440 57458
rect 161388 57394 161440 57400
rect 161400 6914 161428 57394
rect 161308 6886 161428 6914
rect 160376 4004 160428 4010
rect 160376 3946 160428 3952
rect 160192 2848 160244 2854
rect 160192 2790 160244 2796
rect 161308 480 161336 6886
rect 161584 3505 161612 59758
rect 162124 57520 162176 57526
rect 162124 57462 162176 57468
rect 162136 5098 162164 57462
rect 162492 6588 162544 6594
rect 162492 6530 162544 6536
rect 162124 5092 162176 5098
rect 162124 5034 162176 5040
rect 161570 3496 161626 3505
rect 161570 3431 161626 3440
rect 162504 480 162532 6530
rect 162964 3641 162992 59774
rect 163148 59758 163214 59786
rect 164074 59832 164126 59838
rect 164074 59774 164126 59780
rect 164986 59786 165014 60044
rect 165886 59786 165914 60044
rect 166786 59786 166814 60044
rect 167686 59786 167714 60044
rect 164986 59758 165016 59786
rect 163148 57322 163176 59758
rect 164988 57390 165016 59758
rect 165724 59758 165914 59786
rect 166736 59758 166814 59786
rect 167656 59758 167714 59786
rect 168380 59832 168432 59838
rect 168606 59786 168634 60044
rect 169506 59838 169534 60044
rect 168380 59774 168432 59780
rect 164976 57384 165028 57390
rect 164976 57326 165028 57332
rect 163136 57316 163188 57322
rect 163136 57258 163188 57264
rect 165528 57316 165580 57322
rect 165528 57258 165580 57264
rect 164148 10464 164200 10470
rect 164148 10406 164200 10412
rect 162950 3632 163006 3641
rect 162950 3567 163006 3576
rect 164160 3398 164188 10406
rect 165540 3398 165568 57258
rect 163688 3392 163740 3398
rect 163688 3334 163740 3340
rect 164148 3392 164200 3398
rect 164148 3334 164200 3340
rect 164884 3392 164936 3398
rect 164884 3334 164936 3340
rect 165528 3392 165580 3398
rect 165724 3369 165752 59758
rect 166264 57656 166316 57662
rect 166264 57598 166316 57604
rect 166080 6656 166132 6662
rect 166080 6598 166132 6604
rect 165528 3334 165580 3340
rect 165710 3360 165766 3369
rect 163700 480 163728 3334
rect 164896 480 164924 3334
rect 165710 3295 165766 3304
rect 166092 480 166120 6598
rect 166276 6186 166304 57598
rect 166736 57254 166764 59758
rect 167656 57662 167684 59758
rect 167644 57656 167696 57662
rect 167644 57598 167696 57604
rect 166724 57248 166776 57254
rect 166724 57190 166776 57196
rect 168288 10532 168340 10538
rect 168288 10474 168340 10480
rect 166264 6180 166316 6186
rect 166264 6122 166316 6128
rect 168300 3398 168328 10474
rect 168392 4894 168420 59774
rect 168484 59758 168634 59786
rect 169494 59832 169546 59838
rect 170406 59786 170434 60044
rect 169494 59774 169546 59780
rect 169772 59758 170434 59786
rect 171306 59786 171334 60044
rect 172206 59786 172234 60044
rect 173106 59786 173134 60044
rect 171306 59758 171364 59786
rect 168380 4888 168432 4894
rect 168380 4830 168432 4836
rect 168484 4826 168512 59758
rect 169576 14884 169628 14890
rect 169576 14826 169628 14832
rect 168472 4820 168524 4826
rect 168472 4762 168524 4768
rect 168380 4004 168432 4010
rect 168380 3946 168432 3952
rect 167184 3392 167236 3398
rect 167184 3334 167236 3340
rect 168288 3392 168340 3398
rect 168288 3334 168340 3340
rect 167196 480 167224 3334
rect 168392 480 168420 3946
rect 169588 480 169616 14826
rect 169772 4962 169800 59758
rect 171336 57526 171364 59758
rect 172164 59758 172234 59786
rect 172532 59758 173134 59786
rect 173900 59832 173952 59838
rect 174006 59786 174034 60044
rect 174926 59838 174954 60044
rect 173900 59774 173952 59780
rect 171324 57520 171376 57526
rect 171324 57462 171376 57468
rect 172164 56642 172192 59758
rect 170404 56636 170456 56642
rect 170404 56578 170456 56584
rect 172152 56636 172204 56642
rect 172152 56578 172204 56584
rect 170416 28286 170444 56578
rect 170404 28280 170456 28286
rect 170404 28222 170456 28228
rect 170772 10600 170824 10606
rect 170772 10542 170824 10548
rect 169760 4956 169812 4962
rect 169760 4898 169812 4904
rect 170784 480 170812 10542
rect 172532 5030 172560 59758
rect 173808 26920 173860 26926
rect 173808 26862 173860 26868
rect 172520 5024 172572 5030
rect 172520 4966 172572 4972
rect 173820 3398 173848 26862
rect 173912 3874 173940 59774
rect 174004 59758 174034 59786
rect 174914 59832 174966 59838
rect 175826 59786 175854 60044
rect 176726 59786 176754 60044
rect 177626 59786 177654 60044
rect 178526 59786 178554 60044
rect 174914 59774 174966 59780
rect 175292 59758 175854 59786
rect 176672 59758 176754 59786
rect 177592 59758 177654 59786
rect 178052 59758 178554 59786
rect 179426 59786 179454 60044
rect 180346 59786 180374 60044
rect 179426 59758 179460 59786
rect 173900 3868 173952 3874
rect 173900 3810 173952 3816
rect 174004 3806 174032 59758
rect 175188 10668 175240 10674
rect 175188 10610 175240 10616
rect 173992 3800 174044 3806
rect 173992 3742 174044 3748
rect 175200 3398 175228 10610
rect 175292 3942 175320 59758
rect 176672 57458 176700 59758
rect 176660 57452 176712 57458
rect 176660 57394 176712 57400
rect 177304 57452 177356 57458
rect 177304 57394 177356 57400
rect 175280 3936 175332 3942
rect 175280 3878 175332 3884
rect 173164 3392 173216 3398
rect 173164 3334 173216 3340
rect 173808 3392 173860 3398
rect 173808 3334 173860 3340
rect 174268 3392 174320 3398
rect 174268 3334 174320 3340
rect 175188 3392 175240 3398
rect 175188 3334 175240 3340
rect 171968 3256 172020 3262
rect 171968 3198 172020 3204
rect 171980 480 172008 3198
rect 173176 480 173204 3334
rect 174280 480 174308 3334
rect 175464 3324 175516 3330
rect 175464 3266 175516 3272
rect 175476 480 175504 3266
rect 177316 3262 177344 57394
rect 177592 57322 177620 59758
rect 177580 57316 177632 57322
rect 177580 57258 177632 57264
rect 177856 10736 177908 10742
rect 177856 10678 177908 10684
rect 177304 3256 177356 3262
rect 177304 3198 177356 3204
rect 176660 3120 176712 3126
rect 176660 3062 176712 3068
rect 176672 480 176700 3062
rect 177868 480 177896 10678
rect 178052 4010 178080 59758
rect 179432 57458 179460 59758
rect 179524 59758 180374 59786
rect 181246 59786 181274 60044
rect 182146 59786 182174 60044
rect 183046 59786 183074 60044
rect 183946 59786 183974 60044
rect 181246 59758 181300 59786
rect 182146 59758 182220 59786
rect 179420 57452 179472 57458
rect 179420 57394 179472 57400
rect 179328 56636 179380 56642
rect 179328 56578 179380 56584
rect 179340 6914 179368 56578
rect 179064 6886 179368 6914
rect 178040 4004 178092 4010
rect 178040 3946 178092 3952
rect 179064 480 179092 6886
rect 179524 3330 179552 59758
rect 181272 56642 181300 59758
rect 181260 56636 181312 56642
rect 181260 56578 181312 56584
rect 180064 16176 180116 16182
rect 180064 16118 180116 16124
rect 179512 3324 179564 3330
rect 179512 3266 179564 3272
rect 180076 3126 180104 16118
rect 180708 13456 180760 13462
rect 180708 13398 180760 13404
rect 180720 3398 180748 13398
rect 182088 10804 182140 10810
rect 182088 10746 182140 10752
rect 182100 3398 182128 10746
rect 180248 3392 180300 3398
rect 180248 3334 180300 3340
rect 180708 3392 180760 3398
rect 180708 3334 180760 3340
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 182088 3392 182140 3398
rect 182088 3334 182140 3340
rect 180064 3120 180116 3126
rect 180064 3062 180116 3068
rect 180260 480 180288 3334
rect 181456 480 181484 3334
rect 182192 490 182220 59758
rect 183020 59758 183074 59786
rect 183940 59758 183974 59786
rect 184846 59786 184874 60044
rect 185746 59786 185774 60044
rect 186666 59786 186694 60044
rect 187566 59786 187594 60044
rect 188466 59786 188494 60044
rect 184846 59758 184888 59786
rect 185746 59758 185808 59786
rect 186666 59758 186728 59786
rect 187566 59758 187648 59786
rect 183020 57526 183048 59758
rect 183008 57520 183060 57526
rect 183008 57462 183060 57468
rect 183940 57254 183968 59758
rect 184204 57520 184256 57526
rect 184204 57462 184256 57468
rect 183928 57248 183980 57254
rect 183928 57190 183980 57196
rect 184216 3330 184244 57462
rect 184860 4962 184888 59758
rect 185780 57662 185808 59758
rect 185768 57656 185820 57662
rect 185768 57598 185820 57604
rect 186700 56778 186728 59758
rect 186964 57656 187016 57662
rect 186964 57598 187016 57604
rect 186688 56772 186740 56778
rect 186688 56714 186740 56720
rect 186228 10872 186280 10878
rect 186228 10814 186280 10820
rect 184848 4956 184900 4962
rect 184848 4898 184900 4904
rect 186240 3398 186268 10814
rect 186976 6186 187004 57598
rect 187332 6724 187384 6730
rect 187332 6666 187384 6672
rect 186964 6180 187016 6186
rect 186964 6122 187016 6128
rect 184940 3392 184992 3398
rect 184940 3334 184992 3340
rect 186228 3392 186280 3398
rect 186228 3334 186280 3340
rect 184204 3324 184256 3330
rect 184204 3266 184256 3272
rect 183744 3188 183796 3194
rect 183744 3130 183796 3136
rect 182376 598 182588 626
rect 182376 490 182404 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 462 182404 490
rect 182560 480 182588 598
rect 183756 480 183784 3130
rect 184952 480 184980 3334
rect 186136 3324 186188 3330
rect 186136 3266 186188 3272
rect 186148 480 186176 3266
rect 187344 480 187372 6666
rect 187620 4826 187648 59758
rect 188448 59758 188494 59786
rect 189366 59786 189394 60044
rect 190266 59786 190294 60044
rect 191166 59786 191194 60044
rect 192066 59786 192094 60044
rect 189366 59758 189396 59786
rect 190266 59758 190316 59786
rect 191166 59758 191236 59786
rect 188448 57390 188476 59758
rect 188436 57384 188488 57390
rect 188436 57326 188488 57332
rect 189368 57254 189396 59758
rect 190288 57322 190316 59758
rect 191208 57662 191236 59758
rect 192036 59758 192094 59786
rect 192986 59786 193014 60044
rect 193886 59786 193914 60044
rect 192986 59758 193168 59786
rect 192036 57662 192064 59758
rect 191196 57656 191248 57662
rect 191196 57598 191248 57604
rect 191748 57656 191800 57662
rect 191748 57598 191800 57604
rect 192024 57656 192076 57662
rect 192024 57598 192076 57604
rect 193036 57656 193088 57662
rect 193036 57598 193088 57604
rect 190276 57316 190328 57322
rect 190276 57258 190328 57264
rect 188436 57248 188488 57254
rect 188436 57190 188488 57196
rect 189356 57248 189408 57254
rect 189356 57190 189408 57196
rect 188344 56228 188396 56234
rect 188344 56170 188396 56176
rect 187608 4820 187660 4826
rect 187608 4762 187660 4768
rect 188356 3194 188384 56170
rect 188448 4214 188476 57190
rect 191104 56772 191156 56778
rect 191104 56714 191156 56720
rect 188988 10940 189040 10946
rect 188988 10882 189040 10888
rect 188436 4208 188488 4214
rect 188436 4150 188488 4156
rect 189000 3398 189028 10882
rect 191116 4894 191144 56714
rect 191104 4888 191156 4894
rect 191104 4830 191156 4836
rect 191760 4282 191788 57598
rect 192944 11008 192996 11014
rect 192944 10950 192996 10956
rect 191748 4276 191800 4282
rect 191748 4218 191800 4224
rect 189724 4208 189776 4214
rect 189724 4150 189776 4156
rect 188528 3392 188580 3398
rect 188528 3334 188580 3340
rect 188988 3392 189040 3398
rect 188988 3334 189040 3340
rect 188344 3188 188396 3194
rect 188344 3130 188396 3136
rect 188540 480 188568 3334
rect 189736 480 189764 4150
rect 190828 3800 190880 3806
rect 190828 3742 190880 3748
rect 190840 480 190868 3742
rect 192956 3398 192984 10950
rect 193048 4350 193076 57598
rect 193140 4418 193168 59758
rect 193876 59758 193914 59786
rect 194786 59786 194814 60044
rect 195686 59786 195714 60044
rect 196586 59786 196614 60044
rect 197486 59786 197514 60044
rect 194786 59758 194824 59786
rect 195686 59758 195928 59786
rect 196586 59758 196664 59786
rect 193876 57662 193904 59758
rect 194796 57662 194824 59758
rect 193864 57656 193916 57662
rect 193864 57598 193916 57604
rect 194508 57656 194560 57662
rect 194508 57598 194560 57604
rect 194784 57656 194836 57662
rect 194784 57598 194836 57604
rect 195796 57656 195848 57662
rect 195796 57598 195848 57604
rect 194416 9104 194468 9110
rect 194416 9046 194468 9052
rect 193220 4956 193272 4962
rect 193220 4898 193272 4904
rect 193128 4412 193180 4418
rect 193128 4354 193180 4360
rect 193036 4344 193088 4350
rect 193036 4286 193088 4292
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 192944 3392 192996 3398
rect 192944 3334 192996 3340
rect 192036 480 192064 3334
rect 193232 480 193260 4898
rect 194428 480 194456 9046
rect 194520 4486 194548 57598
rect 195612 10260 195664 10266
rect 195612 10202 195664 10208
rect 194508 4480 194560 4486
rect 194508 4422 194560 4428
rect 195624 480 195652 10202
rect 195808 4554 195836 57598
rect 195900 4622 195928 59758
rect 196636 57662 196664 59758
rect 197464 59758 197514 59786
rect 198406 59786 198434 60044
rect 199306 59786 199334 60044
rect 198406 59758 198596 59786
rect 197464 57662 197492 59758
rect 196624 57656 196676 57662
rect 196624 57598 196676 57604
rect 197268 57656 197320 57662
rect 197268 57598 197320 57604
rect 197452 57656 197504 57662
rect 197452 57598 197504 57604
rect 196624 57384 196676 57390
rect 196624 57326 196676 57332
rect 196636 6254 196664 57326
rect 196624 6248 196676 6254
rect 196624 6190 196676 6196
rect 196808 6180 196860 6186
rect 196808 6122 196860 6128
rect 195888 4616 195940 4622
rect 195888 4558 195940 4564
rect 195796 4548 195848 4554
rect 195796 4490 195848 4496
rect 196820 480 196848 6122
rect 197280 4690 197308 57598
rect 197912 9172 197964 9178
rect 197912 9114 197964 9120
rect 197268 4684 197320 4690
rect 197268 4626 197320 4632
rect 197924 480 197952 9114
rect 198568 5506 198596 59758
rect 199304 59758 199334 59786
rect 200206 59786 200234 60044
rect 201106 59786 201134 60044
rect 202006 59786 202034 60044
rect 202906 59786 202934 60044
rect 200206 59758 200252 59786
rect 201106 59758 201356 59786
rect 202006 59758 202092 59786
rect 199304 57662 199332 59758
rect 200224 57662 200252 59758
rect 198648 57656 198700 57662
rect 198648 57598 198700 57604
rect 199292 57656 199344 57662
rect 199292 57598 199344 57604
rect 200028 57656 200080 57662
rect 200028 57598 200080 57604
rect 200212 57656 200264 57662
rect 200212 57598 200264 57604
rect 198556 5500 198608 5506
rect 198556 5442 198608 5448
rect 198660 4758 198688 57598
rect 199936 10192 199988 10198
rect 199936 10134 199988 10140
rect 198648 4752 198700 4758
rect 198648 4694 198700 4700
rect 199948 3398 199976 10134
rect 200040 5438 200068 57598
rect 200028 5432 200080 5438
rect 200028 5374 200080 5380
rect 201328 5302 201356 59758
rect 202064 57662 202092 59758
rect 202892 59758 202934 59786
rect 203806 59786 203834 60044
rect 204726 59786 204754 60044
rect 205626 59786 205654 60044
rect 206526 59786 206554 60044
rect 207426 59786 207454 60044
rect 208326 59786 208354 60044
rect 203806 59758 204116 59786
rect 204726 59758 204760 59786
rect 205626 59758 205680 59786
rect 206526 59758 206968 59786
rect 202892 57662 202920 59758
rect 201408 57656 201460 57662
rect 201408 57598 201460 57604
rect 202052 57656 202104 57662
rect 202052 57598 202104 57604
rect 202788 57656 202840 57662
rect 202788 57598 202840 57604
rect 202880 57656 202932 57662
rect 202880 57598 202932 57604
rect 201420 5370 201448 57598
rect 202144 57316 202196 57322
rect 202144 57258 202196 57264
rect 202156 13122 202184 57258
rect 202144 13116 202196 13122
rect 202144 13058 202196 13064
rect 202696 10124 202748 10130
rect 202696 10066 202748 10072
rect 201500 9240 201552 9246
rect 201500 9182 201552 9188
rect 201408 5364 201460 5370
rect 201408 5306 201460 5312
rect 201316 5296 201368 5302
rect 201316 5238 201368 5244
rect 200304 4888 200356 4894
rect 200304 4830 200356 4836
rect 199108 3392 199160 3398
rect 199108 3334 199160 3340
rect 199936 3392 199988 3398
rect 199936 3334 199988 3340
rect 199120 480 199148 3334
rect 200316 480 200344 4830
rect 201512 480 201540 9182
rect 202708 480 202736 10066
rect 202800 5234 202828 57598
rect 202788 5228 202840 5234
rect 202788 5170 202840 5176
rect 204088 5098 204116 59758
rect 204732 57662 204760 59758
rect 205652 57662 205680 59758
rect 204168 57656 204220 57662
rect 204168 57598 204220 57604
rect 204720 57656 204772 57662
rect 204720 57598 204772 57604
rect 205548 57656 205600 57662
rect 205548 57598 205600 57604
rect 205640 57656 205692 57662
rect 205640 57598 205692 57604
rect 206836 57656 206888 57662
rect 206836 57598 206888 57604
rect 204180 5166 204208 57598
rect 204904 57248 204956 57254
rect 204904 57190 204956 57196
rect 204916 5574 204944 57190
rect 205088 9308 205140 9314
rect 205088 9250 205140 9256
rect 204904 5568 204956 5574
rect 204904 5510 204956 5516
rect 204168 5160 204220 5166
rect 204168 5102 204220 5108
rect 204076 5092 204128 5098
rect 204076 5034 204128 5040
rect 203892 4820 203944 4826
rect 203892 4762 203944 4768
rect 203904 480 203932 4762
rect 205100 480 205128 9250
rect 205560 5030 205588 57598
rect 206744 10056 206796 10062
rect 206744 9998 206796 10004
rect 205548 5024 205600 5030
rect 205548 4966 205600 4972
rect 206756 3398 206784 9998
rect 206848 4962 206876 57598
rect 206836 4956 206888 4962
rect 206836 4898 206888 4904
rect 206940 4894 206968 59758
rect 207400 59758 207454 59786
rect 208228 59758 208354 59786
rect 209226 59786 209254 60044
rect 210126 59786 210154 60044
rect 211046 59786 211074 60044
rect 211946 59786 211974 60044
rect 212846 59786 212874 60044
rect 209226 59758 209268 59786
rect 210126 59758 210188 59786
rect 211046 59758 211108 59786
rect 211946 59758 212028 59786
rect 207400 57662 207428 59758
rect 207388 57656 207440 57662
rect 207388 57598 207440 57604
rect 208228 57322 208256 59758
rect 209240 57662 209268 59758
rect 208308 57656 208360 57662
rect 208308 57598 208360 57604
rect 209228 57656 209280 57662
rect 209228 57598 209280 57604
rect 209688 57656 209740 57662
rect 209688 57598 209740 57604
rect 208216 57316 208268 57322
rect 208216 57258 208268 57264
rect 207388 6248 207440 6254
rect 207388 6190 207440 6196
rect 206928 4888 206980 4894
rect 206928 4830 206980 4836
rect 206192 3392 206244 3398
rect 206192 3334 206244 3340
rect 206744 3392 206796 3398
rect 206744 3334 206796 3340
rect 206204 480 206232 3334
rect 207400 480 207428 6190
rect 208320 4826 208348 57598
rect 209044 29640 209096 29646
rect 209044 29582 209096 29588
rect 208584 9376 208636 9382
rect 208584 9318 208636 9324
rect 208308 4820 208360 4826
rect 208308 4762 208360 4768
rect 208596 480 208624 9318
rect 209056 3806 209084 29582
rect 209700 12442 209728 57598
rect 210160 57254 210188 59758
rect 210148 57248 210200 57254
rect 210148 57190 210200 57196
rect 211080 16318 211108 59758
rect 212000 57186 212028 59758
rect 212828 59758 212874 59786
rect 213746 59786 213774 60044
rect 214646 59786 214674 60044
rect 215546 59786 215574 60044
rect 216466 59786 216494 60044
rect 217366 59786 217394 60044
rect 218266 59786 218294 60044
rect 213746 59758 213776 59786
rect 214646 59758 214696 59786
rect 215546 59758 215616 59786
rect 216466 59758 216628 59786
rect 212828 57662 212856 59758
rect 213748 57934 213776 59758
rect 213736 57928 213788 57934
rect 213736 57870 213788 57876
rect 214668 57662 214696 59758
rect 215588 57662 215616 59758
rect 212816 57656 212868 57662
rect 212816 57598 212868 57604
rect 213828 57656 213880 57662
rect 213828 57598 213880 57604
rect 214656 57656 214708 57662
rect 214656 57598 214708 57604
rect 215208 57656 215260 57662
rect 215208 57598 215260 57604
rect 215576 57656 215628 57662
rect 215576 57598 215628 57604
rect 216496 57656 216548 57662
rect 216496 57598 216548 57604
rect 211988 57180 212040 57186
rect 211988 57122 212040 57128
rect 211068 16312 211120 16318
rect 211068 16254 211120 16260
rect 209688 12436 209740 12442
rect 209688 12378 209740 12384
rect 213840 12374 213868 57598
rect 214472 13116 214524 13122
rect 214472 13058 214524 13064
rect 213828 12368 213880 12374
rect 213828 12310 213880 12316
rect 211068 9988 211120 9994
rect 211068 9930 211120 9936
rect 210976 5568 211028 5574
rect 210976 5510 211028 5516
rect 209044 3800 209096 3806
rect 209044 3742 209096 3748
rect 209780 3392 209832 3398
rect 209780 3334 209832 3340
rect 209792 480 209820 3334
rect 210988 480 211016 5510
rect 211080 3398 211108 9930
rect 213828 9920 213880 9926
rect 213828 9862 213880 9868
rect 212172 9444 212224 9450
rect 212172 9386 212224 9392
rect 211068 3392 211120 3398
rect 211068 3334 211120 3340
rect 212184 480 212212 9386
rect 213840 3398 213868 9862
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 213380 480 213408 3334
rect 214484 480 214512 13058
rect 215220 12306 215248 57598
rect 216508 17474 216536 57598
rect 216496 17468 216548 17474
rect 216496 17410 216548 17416
rect 216600 13666 216628 59758
rect 217336 59758 217394 59786
rect 218256 59758 218294 59786
rect 219166 59786 219194 60044
rect 220066 59786 220094 60044
rect 220966 59786 220994 60044
rect 221866 59786 221894 60044
rect 222786 59786 222814 60044
rect 223686 59786 223714 60044
rect 219166 59758 219204 59786
rect 220066 59758 220124 59786
rect 220966 59758 221044 59786
rect 217336 57662 217364 59758
rect 217324 57656 217376 57662
rect 217324 57598 217376 57604
rect 217968 57656 218020 57662
rect 217968 57598 218020 57604
rect 216588 13660 216640 13666
rect 216588 13602 216640 13608
rect 215208 12300 215260 12306
rect 215208 12242 215260 12248
rect 217980 12170 218008 57598
rect 218256 56642 218284 59758
rect 219176 57458 219204 59758
rect 220096 57662 220124 59758
rect 220084 57656 220136 57662
rect 220084 57598 220136 57604
rect 220728 57656 220780 57662
rect 220728 57598 220780 57604
rect 219164 57452 219216 57458
rect 219164 57394 219216 57400
rect 218244 56636 218296 56642
rect 218244 56578 218296 56584
rect 220084 56636 220136 56642
rect 220084 56578 220136 56584
rect 220096 18698 220124 56578
rect 220084 18692 220136 18698
rect 220084 18634 220136 18640
rect 220636 18624 220688 18630
rect 220636 18566 220688 18572
rect 220084 15972 220136 15978
rect 220084 15914 220136 15920
rect 217968 12164 218020 12170
rect 217968 12106 218020 12112
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 215668 9512 215720 9518
rect 215668 9454 215720 9460
rect 215680 480 215708 9454
rect 218060 4276 218112 4282
rect 218060 4218 218112 4224
rect 216864 4004 216916 4010
rect 216864 3946 216916 3952
rect 216876 480 216904 3946
rect 218072 480 218100 4218
rect 219268 480 219296 9522
rect 220096 4010 220124 15914
rect 220648 6914 220676 18566
rect 220740 13598 220768 57598
rect 221016 56778 221044 59758
rect 221844 59758 221894 59786
rect 222764 59758 222814 59786
rect 223684 59758 223714 59786
rect 224586 59786 224614 60044
rect 225486 59786 225514 60044
rect 226386 59786 226414 60044
rect 227286 59786 227314 60044
rect 228186 59786 228214 60044
rect 229106 59786 229134 60044
rect 230006 59786 230034 60044
rect 230906 59786 230934 60044
rect 231806 59786 231834 60044
rect 232706 59786 232734 60044
rect 224586 59758 224908 59786
rect 225486 59758 225552 59786
rect 226386 59758 226472 59786
rect 227286 59758 227668 59786
rect 228186 59758 228220 59786
rect 229106 59758 229140 59786
rect 230006 59758 230428 59786
rect 230906 59758 230980 59786
rect 221844 57866 221872 59758
rect 221832 57860 221884 57866
rect 221832 57802 221884 57808
rect 222764 57662 222792 59758
rect 223684 57662 223712 59758
rect 222752 57656 222804 57662
rect 222752 57598 222804 57604
rect 223488 57656 223540 57662
rect 223488 57598 223540 57604
rect 223672 57656 223724 57662
rect 223672 57598 223724 57604
rect 224776 57656 224828 57662
rect 224776 57598 224828 57604
rect 222844 57452 222896 57458
rect 222844 57394 222896 57400
rect 221004 56772 221056 56778
rect 221004 56714 221056 56720
rect 222856 25566 222884 57394
rect 222844 25560 222896 25566
rect 222844 25502 222896 25508
rect 220728 13592 220780 13598
rect 220728 13534 220780 13540
rect 223500 12238 223528 57598
rect 224788 21486 224816 57598
rect 224776 21480 224828 21486
rect 224776 21422 224828 21428
rect 224776 19984 224828 19990
rect 224776 19926 224828 19932
rect 223488 12232 223540 12238
rect 223488 12174 223540 12180
rect 222752 9648 222804 9654
rect 222752 9590 222804 9596
rect 220464 6886 220676 6914
rect 220084 4004 220136 4010
rect 220084 3946 220136 3952
rect 220464 480 220492 6886
rect 221556 4344 221608 4350
rect 221556 4286 221608 4292
rect 221568 480 221596 4286
rect 222764 480 222792 9590
rect 224788 2990 224816 19926
rect 224880 13530 224908 59758
rect 225524 57798 225552 59758
rect 225512 57792 225564 57798
rect 225512 57734 225564 57740
rect 226444 57662 226472 59758
rect 226432 57656 226484 57662
rect 226432 57598 226484 57604
rect 227536 57656 227588 57662
rect 227536 57598 227588 57604
rect 224868 13524 224920 13530
rect 224868 13466 224920 13472
rect 227548 13394 227576 57598
rect 227536 13388 227588 13394
rect 227536 13330 227588 13336
rect 227640 12102 227668 59758
rect 228192 57662 228220 59758
rect 229112 57662 229140 59758
rect 228180 57656 228232 57662
rect 228180 57598 228232 57604
rect 229008 57656 229060 57662
rect 229008 57598 229060 57604
rect 229100 57656 229152 57662
rect 229100 57598 229152 57604
rect 230296 57656 230348 57662
rect 230296 57598 230348 57604
rect 228364 56772 228416 56778
rect 228364 56714 228416 56720
rect 228376 20058 228404 56714
rect 228364 20052 228416 20058
rect 228364 19994 228416 20000
rect 227628 12096 227680 12102
rect 227628 12038 227680 12044
rect 226340 8900 226392 8906
rect 226340 8842 226392 8848
rect 225144 4412 225196 4418
rect 225144 4354 225196 4360
rect 223948 2984 224000 2990
rect 223948 2926 224000 2932
rect 224776 2984 224828 2990
rect 224776 2926 224828 2932
rect 223960 480 223988 2926
rect 225156 480 225184 4354
rect 226352 480 226380 8842
rect 229020 6526 229048 57598
rect 229836 8832 229888 8838
rect 229836 8774 229888 8780
rect 229008 6520 229060 6526
rect 229008 6462 229060 6468
rect 228732 4480 228784 4486
rect 228732 4422 228784 4428
rect 227536 3868 227588 3874
rect 227536 3810 227588 3816
rect 227548 480 227576 3810
rect 228744 480 228772 4422
rect 229848 480 229876 8774
rect 230308 6458 230336 57598
rect 230296 6452 230348 6458
rect 230296 6394 230348 6400
rect 230400 6390 230428 59758
rect 230952 57662 230980 59758
rect 231780 59758 231834 59786
rect 232700 59758 232734 59786
rect 233606 59786 233634 60044
rect 234526 59786 234554 60044
rect 235426 59786 235454 60044
rect 236326 59786 236354 60044
rect 237226 59786 237254 60044
rect 233606 59758 233648 59786
rect 234526 59758 234568 59786
rect 235426 59758 235488 59786
rect 236326 59758 236408 59786
rect 230940 57656 230992 57662
rect 230940 57598 230992 57604
rect 231676 57656 231728 57662
rect 231676 57598 231728 57604
rect 230388 6384 230440 6390
rect 230388 6326 230440 6332
rect 231688 6322 231716 57598
rect 231676 6316 231728 6322
rect 231676 6258 231728 6264
rect 231780 6254 231808 59758
rect 232700 57662 232728 59758
rect 232688 57656 232740 57662
rect 232688 57598 232740 57604
rect 233148 57656 233200 57662
rect 233148 57598 233200 57604
rect 231768 6248 231820 6254
rect 231768 6190 231820 6196
rect 233160 6186 233188 57598
rect 233620 57390 233648 59758
rect 233608 57384 233660 57390
rect 233608 57326 233660 57332
rect 233884 33788 233936 33794
rect 233884 33730 233936 33736
rect 233424 8764 233476 8770
rect 233424 8706 233476 8712
rect 233148 6180 233200 6186
rect 233148 6122 233200 6128
rect 232228 4548 232280 4554
rect 232228 4490 232280 4496
rect 231032 3120 231084 3126
rect 231032 3062 231084 3068
rect 231044 480 231072 3062
rect 232240 480 232268 4490
rect 233436 480 233464 8706
rect 233896 3126 233924 33730
rect 234540 13258 234568 59758
rect 235460 57526 235488 59758
rect 236380 57662 236408 59758
rect 237208 59758 237254 59786
rect 238126 59786 238154 60044
rect 239026 59786 239054 60044
rect 239926 59786 239954 60044
rect 240846 59786 240874 60044
rect 241746 59786 241774 60044
rect 238126 59758 238156 59786
rect 239026 59758 239076 59786
rect 239926 59758 239996 59786
rect 240846 59758 240916 59786
rect 236368 57656 236420 57662
rect 236368 57598 236420 57604
rect 235448 57520 235500 57526
rect 235448 57462 235500 57468
rect 237208 56710 237236 59758
rect 238024 57656 238076 57662
rect 238024 57598 238076 57604
rect 237196 56704 237248 56710
rect 237196 56646 237248 56652
rect 238036 22778 238064 57598
rect 238128 57458 238156 59758
rect 238116 57452 238168 57458
rect 238116 57394 238168 57400
rect 238668 57452 238720 57458
rect 238668 57394 238720 57400
rect 238024 22772 238076 22778
rect 238024 22714 238076 22720
rect 238024 21412 238076 21418
rect 238024 21354 238076 21360
rect 234528 13252 234580 13258
rect 234528 13194 234580 13200
rect 237012 8696 237064 8702
rect 237012 8638 237064 8644
rect 235816 4616 235868 4622
rect 235816 4558 235868 4564
rect 234620 4140 234672 4146
rect 234620 4082 234672 4088
rect 233884 3120 233936 3126
rect 233884 3062 233936 3068
rect 234632 480 234660 4082
rect 235828 480 235856 4558
rect 237024 480 237052 8638
rect 238036 3874 238064 21354
rect 238680 11966 238708 57394
rect 239048 57050 239076 59758
rect 239968 57390 239996 59758
rect 240888 57458 240916 59758
rect 241716 59758 241774 59786
rect 242646 59786 242674 60044
rect 243546 59786 243574 60044
rect 244446 59786 244474 60044
rect 245346 59786 245374 60044
rect 246246 59786 246274 60044
rect 247166 59786 247194 60044
rect 242646 59758 242756 59786
rect 243546 59758 243584 59786
rect 244446 59758 244504 59786
rect 245346 59758 245608 59786
rect 241716 57458 241744 59758
rect 240876 57452 240928 57458
rect 240876 57394 240928 57400
rect 241428 57452 241480 57458
rect 241428 57394 241480 57400
rect 241704 57452 241756 57458
rect 241704 57394 241756 57400
rect 239956 57384 240008 57390
rect 239956 57326 240008 57332
rect 239036 57044 239088 57050
rect 239036 56986 239088 56992
rect 240784 56704 240836 56710
rect 240784 56646 240836 56652
rect 240796 14686 240824 56646
rect 241440 24138 241468 57394
rect 241428 24132 241480 24138
rect 241428 24074 241480 24080
rect 240876 16040 240928 16046
rect 240876 15982 240928 15988
rect 240784 14680 240836 14686
rect 240784 14622 240836 14628
rect 238668 11960 238720 11966
rect 238668 11902 238720 11908
rect 240508 8628 240560 8634
rect 240508 8570 240560 8576
rect 239312 4684 239364 4690
rect 239312 4626 239364 4632
rect 238024 3868 238076 3874
rect 238024 3810 238076 3816
rect 238116 3800 238168 3806
rect 238116 3742 238168 3748
rect 238128 480 238156 3742
rect 239324 480 239352 4626
rect 240520 480 240548 8570
rect 240888 4146 240916 15982
rect 242728 7206 242756 59758
rect 243556 57458 243584 59758
rect 244476 57458 244504 59758
rect 242808 57452 242860 57458
rect 242808 57394 242860 57400
rect 243544 57452 243596 57458
rect 243544 57394 243596 57400
rect 244188 57452 244240 57458
rect 244188 57394 244240 57400
rect 244464 57452 244516 57458
rect 244464 57394 244516 57400
rect 245476 57452 245528 57458
rect 245476 57394 245528 57400
rect 242716 7200 242768 7206
rect 242716 7142 242768 7148
rect 242820 7138 242848 57394
rect 244096 8560 244148 8566
rect 244096 8502 244148 8508
rect 242808 7132 242860 7138
rect 242808 7074 242860 7080
rect 242900 4752 242952 4758
rect 242900 4694 242952 4700
rect 240876 4140 240928 4146
rect 240876 4082 240928 4088
rect 241704 3868 241756 3874
rect 241704 3810 241756 3816
rect 241716 480 241744 3810
rect 242912 480 242940 4694
rect 244108 480 244136 8502
rect 244200 7274 244228 57394
rect 245488 7342 245516 57394
rect 245580 7410 245608 59758
rect 246224 59758 246274 59786
rect 247144 59758 247194 59786
rect 248066 59786 248094 60044
rect 248966 59786 248994 60044
rect 249866 59786 249894 60044
rect 250766 59786 250794 60044
rect 251666 59786 251694 60044
rect 252586 59786 252614 60044
rect 248066 59758 248276 59786
rect 248966 59758 249012 59786
rect 249866 59758 249932 59786
rect 250766 59758 251128 59786
rect 246224 57458 246252 59758
rect 246212 57452 246264 57458
rect 246212 57394 246264 57400
rect 246948 57452 247000 57458
rect 246948 57394 247000 57400
rect 246304 57044 246356 57050
rect 246304 56986 246356 56992
rect 246316 14618 246344 56986
rect 246304 14612 246356 14618
rect 246304 14554 246356 14560
rect 246396 14544 246448 14550
rect 246396 14486 246448 14492
rect 245568 7404 245620 7410
rect 245568 7346 245620 7352
rect 245476 7336 245528 7342
rect 245476 7278 245528 7284
rect 244188 7268 244240 7274
rect 244188 7210 244240 7216
rect 246304 5500 246356 5506
rect 246304 5442 246356 5448
rect 245200 3392 245252 3398
rect 245200 3334 245252 3340
rect 245212 480 245240 3334
rect 246316 2802 246344 5442
rect 246408 3398 246436 14486
rect 246960 7478 246988 57394
rect 247144 57390 247172 59758
rect 247132 57384 247184 57390
rect 247132 57326 247184 57332
rect 247592 8492 247644 8498
rect 247592 8434 247644 8440
rect 246948 7472 247000 7478
rect 246948 7414 247000 7420
rect 246396 3392 246448 3398
rect 246396 3334 246448 3340
rect 246316 2774 246436 2802
rect 246408 480 246436 2774
rect 247604 480 247632 8434
rect 248248 8294 248276 59758
rect 248984 57390 249012 59758
rect 249904 57390 249932 59758
rect 248328 57384 248380 57390
rect 248328 57326 248380 57332
rect 248972 57384 249024 57390
rect 248972 57326 249024 57332
rect 249708 57384 249760 57390
rect 249708 57326 249760 57332
rect 249892 57384 249944 57390
rect 249892 57326 249944 57332
rect 250996 57384 251048 57390
rect 250996 57326 251048 57332
rect 248236 8288 248288 8294
rect 248236 8230 248288 8236
rect 248340 7546 248368 57326
rect 249064 56024 249116 56030
rect 249064 55966 249116 55972
rect 248328 7540 248380 7546
rect 248328 7482 248380 7488
rect 249076 3806 249104 55966
rect 249720 8226 249748 57326
rect 249708 8220 249760 8226
rect 249708 8162 249760 8168
rect 251008 8158 251036 57326
rect 250996 8152 251048 8158
rect 250996 8094 251048 8100
rect 251100 8090 251128 59758
rect 251652 59758 251694 59786
rect 252572 59758 252614 59786
rect 253486 59786 253514 60044
rect 254386 59786 254414 60044
rect 255286 59786 255314 60044
rect 256186 59786 256214 60044
rect 257086 59786 257114 60044
rect 253486 59758 253888 59786
rect 254386 59758 254440 59786
rect 255286 59758 255360 59786
rect 256186 59758 256556 59786
rect 251652 57390 251680 59758
rect 252572 57390 252600 59758
rect 251640 57384 251692 57390
rect 251640 57326 251692 57332
rect 252468 57384 252520 57390
rect 252468 57326 252520 57332
rect 252560 57384 252612 57390
rect 252560 57326 252612 57332
rect 253756 57384 253808 57390
rect 253756 57326 253808 57332
rect 251824 54528 251876 54534
rect 251824 54470 251876 54476
rect 251180 8424 251232 8430
rect 251180 8366 251232 8372
rect 251088 8084 251140 8090
rect 251088 8026 251140 8032
rect 249984 5432 250036 5438
rect 249984 5374 250036 5380
rect 249064 3800 249116 3806
rect 249064 3742 249116 3748
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 248800 480 248828 2994
rect 249996 480 250024 5374
rect 251192 480 251220 8366
rect 251836 3058 251864 54470
rect 252480 8022 252508 57326
rect 252468 8016 252520 8022
rect 252468 7958 252520 7964
rect 253768 7954 253796 57326
rect 253756 7948 253808 7954
rect 253756 7890 253808 7896
rect 253860 7886 253888 59758
rect 254412 57390 254440 59758
rect 255332 57390 255360 59758
rect 254400 57384 254452 57390
rect 254400 57326 254452 57332
rect 255228 57384 255280 57390
rect 255228 57326 255280 57332
rect 255320 57384 255372 57390
rect 255320 57326 255372 57332
rect 253848 7880 253900 7886
rect 253848 7822 253900 7828
rect 255240 7818 255268 57326
rect 255228 7812 255280 7818
rect 255228 7754 255280 7760
rect 256528 7682 256556 59758
rect 257080 59758 257114 59786
rect 257986 59786 258014 60044
rect 258906 59786 258934 60044
rect 259806 59786 259834 60044
rect 260706 59786 260734 60044
rect 261606 59786 261634 60044
rect 257986 59758 258028 59786
rect 258906 59758 258948 59786
rect 259806 59758 259868 59786
rect 256608 57384 256660 57390
rect 256608 57326 256660 57332
rect 256620 7750 256648 57326
rect 257080 57118 257108 59758
rect 258000 57390 258028 59758
rect 257988 57384 258040 57390
rect 257988 57326 258040 57332
rect 258920 57322 258948 59758
rect 258724 57316 258776 57322
rect 258724 57258 258776 57264
rect 258908 57316 258960 57322
rect 258908 57258 258960 57264
rect 259368 57316 259420 57322
rect 259368 57258 259420 57264
rect 257068 57112 257120 57118
rect 257068 57054 257120 57060
rect 257988 57112 258040 57118
rect 257988 57054 258040 57060
rect 256608 7744 256660 7750
rect 256608 7686 256660 7692
rect 256516 7676 256568 7682
rect 256516 7618 256568 7624
rect 258000 7614 258028 57054
rect 257988 7608 258040 7614
rect 257988 7550 258040 7556
rect 258736 6118 258764 57258
rect 259276 14952 259328 14958
rect 259276 14894 259328 14900
rect 258724 6112 258776 6118
rect 258724 6054 258776 6060
rect 253480 5364 253532 5370
rect 253480 5306 253532 5312
rect 254676 5364 254728 5370
rect 254676 5306 254728 5312
rect 252376 3936 252428 3942
rect 252376 3878 252428 3884
rect 251824 3052 251876 3058
rect 251824 2994 251876 3000
rect 252388 480 252416 3878
rect 253492 480 253520 5306
rect 254688 480 254716 5306
rect 257068 5296 257120 5302
rect 257068 5238 257120 5244
rect 255872 4072 255924 4078
rect 255872 4014 255924 4020
rect 255884 480 255912 4014
rect 257080 480 257108 5238
rect 259288 3398 259316 14894
rect 259380 14482 259408 57258
rect 259840 55894 259868 59758
rect 260668 59758 260734 59786
rect 261588 59758 261634 59786
rect 262506 59786 262534 60044
rect 263406 59786 263434 60044
rect 264306 59786 264334 60044
rect 265226 59786 265254 60044
rect 266126 59786 266154 60044
rect 267026 59786 267054 60044
rect 262506 59758 262536 59786
rect 263406 59758 263456 59786
rect 264306 59758 264376 59786
rect 265226 59758 265296 59786
rect 266126 59758 266308 59786
rect 260104 56092 260156 56098
rect 260104 56034 260156 56040
rect 259828 55888 259880 55894
rect 259828 55830 259880 55836
rect 259368 14476 259420 14482
rect 259368 14418 259420 14424
rect 260116 3874 260144 56034
rect 260668 11898 260696 59758
rect 261588 57322 261616 59758
rect 261576 57316 261628 57322
rect 261576 57258 261628 57264
rect 262508 55962 262536 59758
rect 262864 57112 262916 57118
rect 262864 57054 262916 57060
rect 262496 55956 262548 55962
rect 262496 55898 262548 55904
rect 260656 11892 260708 11898
rect 260656 11834 260708 11840
rect 261760 6860 261812 6866
rect 261760 6802 261812 6808
rect 260656 5228 260708 5234
rect 260656 5170 260708 5176
rect 260104 3868 260156 3874
rect 260104 3810 260156 3816
rect 259460 3800 259512 3806
rect 259460 3742 259512 3748
rect 258264 3392 258316 3398
rect 258264 3334 258316 3340
rect 259276 3392 259328 3398
rect 259276 3334 259328 3340
rect 258276 480 258304 3334
rect 259472 480 259500 3742
rect 260668 480 260696 5170
rect 261772 480 261800 6802
rect 262876 5370 262904 57054
rect 263428 11830 263456 59758
rect 264244 57248 264296 57254
rect 264244 57190 264296 57196
rect 263416 11824 263468 11830
rect 263416 11766 263468 11772
rect 264256 6050 264284 57190
rect 264348 57050 264376 59758
rect 265268 57254 265296 59758
rect 265256 57248 265308 57254
rect 265256 57190 265308 57196
rect 264336 57044 264388 57050
rect 264336 56986 264388 56992
rect 264888 57044 264940 57050
rect 264888 56986 264940 56992
rect 264336 13184 264388 13190
rect 264336 13126 264388 13132
rect 264244 6044 264296 6050
rect 264244 5986 264296 5992
rect 262864 5364 262916 5370
rect 262864 5306 262916 5312
rect 264152 5160 264204 5166
rect 264152 5102 264204 5108
rect 262956 3392 263008 3398
rect 262956 3334 263008 3340
rect 262968 480 262996 3334
rect 264164 480 264192 5102
rect 264348 3398 264376 13126
rect 264900 13122 264928 56986
rect 264888 13116 264940 13122
rect 264888 13058 264940 13064
rect 265348 6792 265400 6798
rect 265348 6734 265400 6740
rect 264336 3392 264388 3398
rect 264336 3334 264388 3340
rect 265360 480 265388 6734
rect 266280 4282 266308 59758
rect 267016 59758 267054 59786
rect 267926 59786 267954 60044
rect 268826 59786 268854 60044
rect 269726 59786 269754 60044
rect 270646 59786 270674 60044
rect 271546 59786 271574 60044
rect 272446 59786 272474 60044
rect 267926 59758 267964 59786
rect 268826 59758 268976 59786
rect 269726 59758 269804 59786
rect 270646 59758 270724 59786
rect 271546 59758 271828 59786
rect 267016 57050 267044 59758
rect 267936 57050 267964 59758
rect 267004 57044 267056 57050
rect 267004 56986 267056 56992
rect 267648 57044 267700 57050
rect 267648 56986 267700 56992
rect 267924 57044 267976 57050
rect 267924 56986 267976 56992
rect 267004 37936 267056 37942
rect 267004 37878 267056 37884
rect 266268 4276 266320 4282
rect 266268 4218 266320 4224
rect 266544 4004 266596 4010
rect 266544 3946 266596 3952
rect 266556 480 266584 3946
rect 267016 3942 267044 37878
rect 267660 4350 267688 56986
rect 268844 13728 268896 13734
rect 268844 13670 268896 13676
rect 267740 5092 267792 5098
rect 267740 5034 267792 5040
rect 267648 4344 267700 4350
rect 267648 4286 267700 4292
rect 267004 3936 267056 3942
rect 267004 3878 267056 3884
rect 267752 480 267780 5034
rect 268856 480 268884 13670
rect 268948 4486 268976 59758
rect 269776 57050 269804 59758
rect 270696 57050 270724 59758
rect 269028 57044 269080 57050
rect 269028 56986 269080 56992
rect 269764 57044 269816 57050
rect 269764 56986 269816 56992
rect 270408 57044 270460 57050
rect 270408 56986 270460 56992
rect 270684 57044 270736 57050
rect 270684 56986 270736 56992
rect 271696 57044 271748 57050
rect 271696 56986 271748 56992
rect 268936 4480 268988 4486
rect 268936 4422 268988 4428
rect 269040 4418 269068 56986
rect 269764 17332 269816 17338
rect 269764 17274 269816 17280
rect 269028 4412 269080 4418
rect 269028 4354 269080 4360
rect 269776 4078 269804 17274
rect 270420 4554 270448 56986
rect 271708 5030 271736 56986
rect 271236 5024 271288 5030
rect 271236 4966 271288 4972
rect 271696 5024 271748 5030
rect 271696 4966 271748 4972
rect 270408 4548 270460 4554
rect 270408 4490 270460 4496
rect 269764 4072 269816 4078
rect 269764 4014 269816 4020
rect 270040 3868 270092 3874
rect 270040 3810 270092 3816
rect 270052 480 270080 3810
rect 271248 480 271276 4966
rect 271800 4622 271828 59758
rect 272444 59758 272474 59786
rect 273346 59786 273374 60044
rect 274246 59786 274274 60044
rect 275146 59786 275174 60044
rect 276046 59786 276074 60044
rect 273346 59758 273392 59786
rect 274246 59758 274588 59786
rect 275146 59758 275232 59786
rect 272444 57050 272472 59758
rect 272432 57044 272484 57050
rect 272432 56986 272484 56992
rect 273168 57044 273220 57050
rect 273168 56986 273220 56992
rect 272616 4888 272668 4894
rect 272616 4830 272668 4836
rect 271788 4616 271840 4622
rect 271788 4558 271840 4564
rect 272628 2530 272656 4830
rect 273180 4690 273208 56986
rect 273364 56642 273392 59758
rect 273352 56636 273404 56642
rect 273352 56578 273404 56584
rect 274456 56636 274508 56642
rect 274456 56578 274508 56584
rect 274468 5506 274496 56578
rect 274456 5500 274508 5506
rect 274456 5442 274508 5448
rect 274560 5438 274588 59758
rect 275204 56642 275232 59758
rect 276032 59758 276074 59786
rect 276966 59786 276994 60044
rect 277866 59786 277894 60044
rect 278766 59786 278794 60044
rect 279666 59786 279694 60044
rect 280566 59786 280594 60044
rect 281466 59786 281494 60044
rect 276966 59758 277256 59786
rect 277866 59758 277900 59786
rect 278766 59758 278820 59786
rect 279666 59758 280016 59786
rect 276032 56642 276060 59758
rect 275192 56636 275244 56642
rect 275192 56578 275244 56584
rect 275928 56636 275980 56642
rect 275928 56578 275980 56584
rect 276020 56636 276072 56642
rect 276020 56578 276072 56584
rect 274548 5432 274600 5438
rect 274548 5374 274600 5380
rect 275940 5370 275968 56578
rect 277124 9852 277176 9858
rect 277124 9794 277176 9800
rect 275928 5364 275980 5370
rect 275928 5306 275980 5312
rect 274824 4956 274876 4962
rect 274824 4898 274876 4904
rect 273168 4684 273220 4690
rect 273168 4626 273220 4632
rect 273628 4072 273680 4078
rect 273628 4014 273680 4020
rect 272444 2502 272656 2530
rect 272444 480 272472 2502
rect 273640 480 273668 4014
rect 274836 480 274864 4898
rect 277136 3398 277164 9794
rect 277228 5234 277256 59758
rect 277872 56642 277900 59758
rect 278136 56976 278188 56982
rect 278136 56918 278188 56924
rect 277308 56636 277360 56642
rect 277308 56578 277360 56584
rect 277860 56636 277912 56642
rect 277860 56578 277912 56584
rect 277320 5302 277348 56578
rect 278148 51074 278176 56918
rect 278792 56642 278820 59758
rect 278688 56636 278740 56642
rect 278688 56578 278740 56584
rect 278780 56636 278832 56642
rect 278780 56578 278832 56584
rect 278056 51046 278176 51074
rect 277308 5296 277360 5302
rect 277308 5238 277360 5244
rect 277216 5228 277268 5234
rect 277216 5170 277268 5176
rect 278056 4894 278084 51046
rect 278044 4888 278096 4894
rect 278044 4830 278096 4836
rect 278320 4752 278372 4758
rect 278320 4694 278372 4700
rect 277216 3936 277268 3942
rect 277216 3878 277268 3884
rect 276020 3392 276072 3398
rect 276020 3334 276072 3340
rect 277124 3392 277176 3398
rect 277124 3334 277176 3340
rect 276032 480 276060 3334
rect 277228 1986 277256 3878
rect 277136 1958 277256 1986
rect 277136 480 277164 1958
rect 278332 480 278360 4694
rect 278700 4214 278728 56578
rect 279516 9784 279568 9790
rect 279516 9726 279568 9732
rect 278688 4208 278740 4214
rect 278688 4150 278740 4156
rect 279528 480 279556 9726
rect 279988 5166 280016 59758
rect 280540 59758 280594 59786
rect 281460 59758 281494 59786
rect 282366 59786 282394 60044
rect 283286 59786 283314 60044
rect 284186 59786 284214 60044
rect 285086 59786 285114 60044
rect 285986 59786 286014 60044
rect 286886 59786 286914 60044
rect 287786 59786 287814 60044
rect 288706 59922 288734 60044
rect 282366 59758 282408 59786
rect 280540 56642 280568 59758
rect 280068 56636 280120 56642
rect 280068 56578 280120 56584
rect 280528 56636 280580 56642
rect 280528 56578 280580 56584
rect 281356 56636 281408 56642
rect 281356 56578 281408 56584
rect 279976 5160 280028 5166
rect 279976 5102 280028 5108
rect 280080 5098 280108 56578
rect 281264 13320 281316 13326
rect 281264 13262 281316 13268
rect 280068 5092 280120 5098
rect 280068 5034 280120 5040
rect 281276 3398 281304 13262
rect 281368 4962 281396 56578
rect 281356 4956 281408 4962
rect 281356 4898 281408 4904
rect 281460 4894 281488 59758
rect 282380 56642 282408 59758
rect 282932 59758 283314 59786
rect 283392 59758 284214 59786
rect 284312 59758 285114 59786
rect 285692 59758 286014 59786
rect 286152 59758 286914 59786
rect 287072 59758 287814 59786
rect 288452 59894 288734 59922
rect 282368 56636 282420 56642
rect 282368 56578 282420 56584
rect 282828 56636 282880 56642
rect 282828 56578 282880 56584
rect 282184 56160 282236 56166
rect 282184 56102 282236 56108
rect 281448 4888 281500 4894
rect 281448 4830 281500 4836
rect 281908 4820 281960 4826
rect 281908 4762 281960 4768
rect 280712 3392 280764 3398
rect 280712 3334 280764 3340
rect 281264 3392 281316 3398
rect 281264 3334 281316 3340
rect 280724 480 280752 3334
rect 281920 480 281948 4762
rect 282196 4010 282224 56102
rect 282840 4826 282868 56578
rect 282932 7070 282960 59758
rect 283392 45554 283420 59758
rect 283024 45526 283420 45554
rect 283024 8974 283052 45526
rect 284312 9042 284340 59758
rect 284944 56908 284996 56914
rect 284944 56850 284996 56856
rect 284300 9036 284352 9042
rect 284300 8978 284352 8984
rect 283012 8968 283064 8974
rect 283012 8910 283064 8916
rect 282920 7064 282972 7070
rect 282920 7006 282972 7012
rect 283104 7064 283156 7070
rect 283104 7006 283156 7012
rect 282828 4820 282880 4826
rect 282828 4762 282880 4768
rect 282184 4004 282236 4010
rect 282184 3946 282236 3952
rect 283116 480 283144 7006
rect 284956 5982 284984 56850
rect 285692 14754 285720 59758
rect 286152 45554 286180 59758
rect 285784 45526 286180 45554
rect 285784 36582 285812 45526
rect 285772 36576 285824 36582
rect 285772 36518 285824 36524
rect 286324 36576 286376 36582
rect 286324 36518 286376 36524
rect 285680 14748 285732 14754
rect 285680 14690 285732 14696
rect 285588 12028 285640 12034
rect 285588 11970 285640 11976
rect 285404 6112 285456 6118
rect 285404 6054 285456 6060
rect 284944 5976 284996 5982
rect 284944 5918 284996 5924
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 284312 480 284340 3130
rect 285416 480 285444 6054
rect 285600 3194 285628 11970
rect 286336 3806 286364 36518
rect 287072 14822 287100 59758
rect 288452 57594 288480 59894
rect 289606 59786 289634 60044
rect 290506 59786 290534 60044
rect 288544 59758 289634 59786
rect 290476 59758 290534 59786
rect 291200 59832 291252 59838
rect 291406 59786 291434 60044
rect 292306 59838 292334 60044
rect 291200 59774 291252 59780
rect 288440 57588 288492 57594
rect 288440 57530 288492 57536
rect 287704 57180 287756 57186
rect 287704 57122 287756 57128
rect 287060 14816 287112 14822
rect 287060 14758 287112 14764
rect 287716 6662 287744 57122
rect 288544 31074 288572 59758
rect 290476 57730 290504 59758
rect 290464 57724 290516 57730
rect 290464 57666 290516 57672
rect 289084 57588 289136 57594
rect 289084 57530 289136 57536
rect 288532 31068 288584 31074
rect 288532 31010 288584 31016
rect 289096 14890 289124 57530
rect 289176 28280 289228 28286
rect 289176 28222 289228 28228
rect 289084 14884 289136 14890
rect 289084 14826 289136 14832
rect 287796 14816 287848 14822
rect 287796 14758 287848 14764
rect 287704 6656 287756 6662
rect 287704 6598 287756 6604
rect 286600 6112 286652 6118
rect 286600 6054 286652 6060
rect 286324 3800 286376 3806
rect 286324 3742 286376 3748
rect 285588 3188 285640 3194
rect 285588 3130 285640 3136
rect 286612 480 286640 6054
rect 287808 4078 287836 14758
rect 288992 12436 289044 12442
rect 288992 12378 289044 12384
rect 287796 4072 287848 4078
rect 287796 4014 287848 4020
rect 287796 3324 287848 3330
rect 287796 3266 287848 3272
rect 287808 480 287836 3266
rect 289004 480 289032 12378
rect 289188 3874 289216 28222
rect 290188 6656 290240 6662
rect 290188 6598 290240 6604
rect 289176 3868 289228 3874
rect 289176 3810 289228 3816
rect 290200 480 290228 6598
rect 291212 6594 291240 59774
rect 291304 59758 291434 59786
rect 292294 59832 292346 59838
rect 292294 59774 292346 59780
rect 293206 59786 293234 60044
rect 294106 59922 294134 60044
rect 293972 59894 294134 59922
rect 293206 59758 293264 59786
rect 291304 32434 291332 59758
rect 293236 57186 293264 59758
rect 293972 57594 294000 59894
rect 295026 59786 295054 60044
rect 295926 59786 295954 60044
rect 296826 59786 296854 60044
rect 294064 59758 295054 59786
rect 295444 59758 295954 59786
rect 296824 59758 296854 59786
rect 297726 59786 297754 60044
rect 298626 59786 298654 60044
rect 297726 59758 297772 59786
rect 293960 57588 294012 57594
rect 293960 57530 294012 57536
rect 293224 57180 293276 57186
rect 293224 57122 293276 57128
rect 291292 32428 291344 32434
rect 291292 32370 291344 32376
rect 294064 26926 294092 59758
rect 294052 26920 294104 26926
rect 294052 26862 294104 26868
rect 294604 17400 294656 17406
rect 294604 17342 294656 17348
rect 291844 16108 291896 16114
rect 291844 16050 291896 16056
rect 291200 6588 291252 6594
rect 291200 6530 291252 6536
rect 291856 3942 291884 16050
rect 292488 14748 292540 14754
rect 292488 14690 292540 14696
rect 291844 3936 291896 3942
rect 291844 3878 291896 3884
rect 292500 3398 292528 14690
rect 293684 6588 293736 6594
rect 293684 6530 293736 6536
rect 292580 6044 292632 6050
rect 292580 5986 292632 5992
rect 291384 3392 291436 3398
rect 291384 3334 291436 3340
rect 292488 3392 292540 3398
rect 292488 3334 292540 3340
rect 291396 480 291424 3334
rect 292592 480 292620 5986
rect 293696 480 293724 6530
rect 294616 3330 294644 17342
rect 295444 16182 295472 59758
rect 296824 56642 296852 59758
rect 295984 56636 296036 56642
rect 295984 56578 296036 56584
rect 296812 56636 296864 56642
rect 296812 56578 296864 56584
rect 295616 16312 295668 16318
rect 295616 16254 295668 16260
rect 295432 16176 295484 16182
rect 295432 16118 295484 16124
rect 294880 3800 294932 3806
rect 294880 3742 294932 3748
rect 294604 3324 294656 3330
rect 294604 3266 294656 3272
rect 294892 480 294920 3742
rect 295628 490 295656 16254
rect 295996 13462 296024 56578
rect 297744 56234 297772 59758
rect 298112 59758 298654 59786
rect 299526 59786 299554 60044
rect 300426 59786 300454 60044
rect 301346 59786 301374 60044
rect 299526 59758 299612 59786
rect 297732 56228 297784 56234
rect 297732 56170 297784 56176
rect 295984 13456 296036 13462
rect 295984 13398 296036 13404
rect 298112 6730 298140 59758
rect 298744 57724 298796 57730
rect 298744 57666 298796 57672
rect 298756 6866 298784 57666
rect 299480 57588 299532 57594
rect 299480 57530 299532 57536
rect 299492 9110 299520 57530
rect 299584 29646 299612 59758
rect 300412 59758 300454 59786
rect 300872 59758 301374 59786
rect 302246 59786 302274 60044
rect 303146 59786 303174 60044
rect 303620 59900 303672 59906
rect 303620 59842 303672 59848
rect 302246 59758 302372 59786
rect 300412 57594 300440 59758
rect 300400 57588 300452 57594
rect 300400 57530 300452 57536
rect 299572 29640 299624 29646
rect 299572 29582 299624 29588
rect 300124 26920 300176 26926
rect 300124 26862 300176 26868
rect 299480 9104 299532 9110
rect 299480 9046 299532 9052
rect 298744 6860 298796 6866
rect 298744 6802 298796 6808
rect 298100 6724 298152 6730
rect 298100 6666 298152 6672
rect 297272 6044 297324 6050
rect 297272 5986 297324 5992
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 5986
rect 299664 5976 299716 5982
rect 299664 5918 299716 5924
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 298480 480 298508 3334
rect 299676 480 299704 5918
rect 300136 3398 300164 26862
rect 300872 9178 300900 59758
rect 302344 9246 302372 59758
rect 302436 59758 303174 59786
rect 302436 9314 302464 59758
rect 303160 12368 303212 12374
rect 303160 12310 303212 12316
rect 302424 9308 302476 9314
rect 302424 9250 302476 9256
rect 302332 9240 302384 9246
rect 302332 9182 302384 9188
rect 300860 9172 300912 9178
rect 300860 9114 300912 9120
rect 300768 6724 300820 6730
rect 300768 6666 300820 6672
rect 300124 3392 300176 3398
rect 300124 3334 300176 3340
rect 300780 480 300808 6666
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 301976 480 302004 3878
rect 303172 480 303200 12310
rect 303632 9450 303660 59842
rect 304046 59786 304074 60044
rect 304946 59906 304974 60044
rect 304934 59900 304986 59906
rect 304934 59842 304986 59848
rect 305846 59786 305874 60044
rect 306766 59786 306794 60044
rect 303724 59758 304074 59786
rect 305012 59758 305874 59786
rect 306392 59758 306794 59786
rect 307666 59786 307694 60044
rect 308566 59786 308594 60044
rect 309466 59786 309494 60044
rect 310366 59786 310394 60044
rect 311266 59786 311294 60044
rect 312166 59786 312194 60044
rect 313086 59786 313114 60044
rect 313986 59786 314014 60044
rect 314886 59786 314914 60044
rect 315786 59786 315814 60044
rect 316686 59786 316714 60044
rect 317586 59922 317614 60044
rect 307666 59758 307708 59786
rect 303620 9444 303672 9450
rect 303620 9386 303672 9392
rect 303724 9382 303752 59758
rect 305012 9518 305040 59758
rect 305644 57928 305696 57934
rect 305644 57870 305696 57876
rect 305000 9512 305052 9518
rect 305000 9454 305052 9460
rect 303712 9376 303764 9382
rect 303712 9318 303764 9324
rect 305656 8362 305684 57870
rect 306392 9586 306420 59758
rect 307680 57730 307708 59758
rect 307772 59758 308594 59786
rect 309244 59758 309494 59786
rect 309612 59758 310394 59786
rect 310532 59758 311294 59786
rect 311912 59758 312194 59786
rect 312280 59758 313114 59786
rect 313292 59758 314014 59786
rect 314764 59758 314914 59786
rect 315776 59758 315814 59786
rect 316052 59758 316714 59786
rect 317432 59894 317614 59922
rect 306472 57724 306524 57730
rect 306472 57666 306524 57672
rect 307668 57724 307720 57730
rect 307668 57666 307720 57672
rect 306484 9654 306512 57666
rect 306472 9648 306524 9654
rect 306472 9590 306524 9596
rect 306380 9580 306432 9586
rect 306380 9522 306432 9528
rect 307772 8906 307800 59758
rect 307760 8900 307812 8906
rect 307760 8842 307812 8848
rect 309244 8838 309272 59758
rect 309612 45554 309640 59758
rect 309336 45526 309640 45554
rect 309232 8832 309284 8838
rect 309232 8774 309284 8780
rect 309336 8770 309364 45526
rect 309784 12300 309836 12306
rect 309784 12242 309836 12248
rect 309324 8764 309376 8770
rect 309324 8706 309376 8712
rect 305644 8356 305696 8362
rect 305644 8298 305696 8304
rect 306748 8356 306800 8362
rect 306748 8298 306800 8304
rect 304356 6860 304408 6866
rect 304356 6802 304408 6808
rect 304368 480 304396 6802
rect 305552 4004 305604 4010
rect 305552 3946 305604 3952
rect 305564 480 305592 3946
rect 306760 480 306788 8298
rect 307944 5976 307996 5982
rect 307944 5918 307996 5924
rect 307956 480 307984 5918
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 309060 480 309088 3810
rect 309796 490 309824 12242
rect 310532 8702 310560 59758
rect 310520 8696 310572 8702
rect 310520 8638 310572 8644
rect 311912 8634 311940 59758
rect 312280 45554 312308 59758
rect 312004 45526 312308 45554
rect 311900 8628 311952 8634
rect 311900 8570 311952 8576
rect 312004 8566 312032 45526
rect 312636 8968 312688 8974
rect 312636 8910 312688 8916
rect 311992 8560 312044 8566
rect 311992 8502 312044 8508
rect 311440 5908 311492 5914
rect 311440 5850 311492 5856
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 5850
rect 312648 480 312676 8910
rect 313292 8498 313320 59758
rect 313372 17468 313424 17474
rect 313372 17410 313424 17416
rect 313384 16574 313412 17410
rect 313384 16546 313872 16574
rect 313280 8492 313332 8498
rect 313280 8434 313332 8440
rect 313844 480 313872 16546
rect 314764 8430 314792 59758
rect 315776 57118 315804 59758
rect 315764 57112 315816 57118
rect 315764 57054 315816 57060
rect 316052 14958 316080 59758
rect 317432 57594 317460 59894
rect 318486 59786 318514 60044
rect 319406 59786 319434 60044
rect 320306 59922 320334 60044
rect 317524 59758 318514 59786
rect 319364 59758 319434 59786
rect 320192 59894 320334 59922
rect 317420 57588 317472 57594
rect 317420 57530 317472 57536
rect 316684 56908 316736 56914
rect 316684 56850 316736 56856
rect 316040 14952 316092 14958
rect 316040 14894 316092 14900
rect 316696 13734 316724 56850
rect 316684 13728 316736 13734
rect 316684 13670 316736 13676
rect 316040 13660 316092 13666
rect 316040 13602 316092 13608
rect 314752 8424 314804 8430
rect 314752 8366 314804 8372
rect 315028 5840 315080 5846
rect 315028 5782 315080 5788
rect 315040 480 315068 5782
rect 316052 3398 316080 13602
rect 316776 13456 316828 13462
rect 316776 13398 316828 13404
rect 316788 4010 316816 13398
rect 317524 6798 317552 59758
rect 319364 56914 319392 59758
rect 320192 57050 320220 59894
rect 321206 59786 321234 60044
rect 322106 59786 322134 60044
rect 320284 59758 321234 59786
rect 321572 59758 322134 59786
rect 323006 59786 323034 60044
rect 323906 59786 323934 60044
rect 324826 59786 324854 60044
rect 323006 59758 323072 59786
rect 320180 57044 320232 57050
rect 320180 56986 320232 56992
rect 319352 56908 319404 56914
rect 319352 56850 319404 56856
rect 318064 54596 318116 54602
rect 318064 54538 318116 54544
rect 317512 6792 317564 6798
rect 317512 6734 317564 6740
rect 316776 4004 316828 4010
rect 316776 3946 316828 3952
rect 318076 3806 318104 54538
rect 320284 9858 320312 59758
rect 320824 31068 320876 31074
rect 320824 31010 320876 31016
rect 320456 12164 320508 12170
rect 320456 12106 320508 12112
rect 320272 9852 320324 9858
rect 320272 9794 320324 9800
rect 318524 6792 318576 6798
rect 318524 6734 318576 6740
rect 318064 3800 318116 3806
rect 318064 3742 318116 3748
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 316224 3188 316276 3194
rect 316224 3130 316276 3136
rect 316236 480 316264 3130
rect 317340 480 317368 3334
rect 318536 480 318564 6734
rect 319720 3392 319772 3398
rect 319720 3334 319772 3340
rect 319732 480 319760 3334
rect 320468 490 320496 12106
rect 320836 3942 320864 31010
rect 321572 9790 321600 59758
rect 322204 57860 322256 57866
rect 322204 57802 322256 57808
rect 321560 9784 321612 9790
rect 321560 9726 321612 9732
rect 322216 9042 322244 57802
rect 322940 57588 322992 57594
rect 322940 57530 322992 57536
rect 322296 12164 322348 12170
rect 322296 12106 322348 12112
rect 322204 9036 322256 9042
rect 322204 8978 322256 8984
rect 322112 5772 322164 5778
rect 322112 5714 322164 5720
rect 320824 3936 320876 3942
rect 320824 3878 320876 3884
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 5714
rect 322308 3194 322336 12106
rect 322952 6118 322980 57530
rect 323044 7070 323072 59758
rect 323872 59758 323934 59786
rect 324332 59758 324854 59786
rect 325726 59786 325754 60044
rect 326626 59786 326654 60044
rect 327526 59786 327554 60044
rect 325726 59758 325832 59786
rect 326626 59758 326660 59786
rect 323872 57594 323900 59758
rect 323860 57588 323912 57594
rect 323860 57530 323912 57536
rect 323584 16176 323636 16182
rect 323584 16118 323636 16124
rect 323032 7064 323084 7070
rect 323032 7006 323084 7012
rect 322940 6112 322992 6118
rect 322940 6054 322992 6060
rect 323308 3800 323360 3806
rect 323308 3742 323360 3748
rect 322296 3188 322348 3194
rect 322296 3130 322348 3136
rect 323320 480 323348 3742
rect 323596 3398 323624 16118
rect 324332 6662 324360 59758
rect 325700 57588 325752 57594
rect 325700 57530 325752 57536
rect 324412 18692 324464 18698
rect 324412 18634 324464 18640
rect 324320 6656 324372 6662
rect 324320 6598 324372 6604
rect 323584 3392 323636 3398
rect 323584 3334 323636 3340
rect 324424 480 324452 18634
rect 325608 9104 325660 9110
rect 325608 9046 325660 9052
rect 325620 480 325648 9046
rect 325712 6050 325740 57530
rect 325804 6594 325832 59758
rect 326632 57594 326660 59758
rect 327092 59758 327554 59786
rect 328426 59786 328454 60044
rect 329326 59786 329354 60044
rect 330226 59786 330254 60044
rect 331146 59786 331174 60044
rect 332046 59786 332074 60044
rect 332946 59786 332974 60044
rect 333846 59786 333874 60044
rect 334746 59786 334774 60044
rect 335646 59786 335674 60044
rect 328426 59758 328500 59786
rect 326620 57588 326672 57594
rect 326620 57530 326672 57536
rect 327092 6730 327120 59758
rect 327172 25560 327224 25566
rect 327172 25502 327224 25508
rect 327184 16574 327212 25502
rect 327184 16546 328040 16574
rect 327080 6724 327132 6730
rect 327080 6666 327132 6672
rect 325792 6588 325844 6594
rect 325792 6530 325844 6536
rect 325700 6044 325752 6050
rect 325700 5986 325752 5992
rect 326804 3392 326856 3398
rect 326804 3334 326856 3340
rect 326816 480 326844 3334
rect 328012 480 328040 16546
rect 328472 6866 328500 59758
rect 328564 59758 329354 59786
rect 329852 59758 330254 59786
rect 331140 59758 331174 59786
rect 331232 59758 332074 59786
rect 332704 59758 332974 59786
rect 333808 59758 333874 59786
rect 333992 59758 334774 59786
rect 335464 59758 335674 59786
rect 336546 59786 336574 60044
rect 337466 59786 337494 60044
rect 338366 59786 338394 60044
rect 339266 59786 339294 60044
rect 340166 59786 340194 60044
rect 336546 59758 336596 59786
rect 337466 59758 337516 59786
rect 338366 59758 338436 59786
rect 339266 59758 339448 59786
rect 328460 6860 328512 6866
rect 328460 6802 328512 6808
rect 328564 5982 328592 59758
rect 328552 5976 328604 5982
rect 328552 5918 328604 5924
rect 329852 5914 329880 59758
rect 331140 57594 331168 59758
rect 329932 57588 329984 57594
rect 329932 57530 329984 57536
rect 331128 57588 331180 57594
rect 331128 57530 331180 57536
rect 329840 5908 329892 5914
rect 329840 5850 329892 5856
rect 329944 5846 329972 57530
rect 331232 6798 331260 59758
rect 331864 57724 331916 57730
rect 331864 57666 331916 57672
rect 331588 13592 331640 13598
rect 331588 13534 331640 13540
rect 331220 6792 331272 6798
rect 331220 6734 331272 6740
rect 329932 5840 329984 5846
rect 329932 5782 329984 5788
rect 329196 5568 329248 5574
rect 329196 5510 329248 5516
rect 329208 480 329236 5510
rect 330392 3936 330444 3942
rect 330392 3878 330444 3884
rect 330404 480 330432 3878
rect 331600 480 331628 13534
rect 331876 9110 331904 57666
rect 331864 9104 331916 9110
rect 331864 9046 331916 9052
rect 332704 5778 332732 59758
rect 333808 57730 333836 59758
rect 333796 57724 333848 57730
rect 333796 57666 333848 57672
rect 332692 5772 332744 5778
rect 332692 5714 332744 5720
rect 332692 5636 332744 5642
rect 332692 5578 332744 5584
rect 332704 480 332732 5578
rect 333992 5574 334020 59758
rect 335360 57588 335412 57594
rect 335360 57530 335412 57536
rect 334072 20052 334124 20058
rect 334072 19994 334124 20000
rect 334084 16574 334112 19994
rect 334084 16546 334664 16574
rect 333980 5568 334032 5574
rect 333980 5510 334032 5516
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 333900 480 333928 3946
rect 334636 490 334664 16546
rect 335372 3482 335400 57530
rect 335464 5642 335492 59758
rect 336568 57594 336596 59758
rect 337488 57594 337516 59758
rect 338408 57594 338436 59758
rect 336556 57588 336608 57594
rect 336556 57530 336608 57536
rect 337476 57588 337528 57594
rect 337476 57530 337528 57536
rect 338028 57588 338080 57594
rect 338028 57530 338080 57536
rect 338396 57588 338448 57594
rect 338396 57530 338448 57536
rect 339316 57588 339368 57594
rect 339316 57530 339368 57536
rect 335452 5636 335504 5642
rect 335452 5578 335504 5584
rect 338040 5574 338068 57530
rect 338672 9036 338724 9042
rect 338672 8978 338724 8984
rect 338028 5568 338080 5574
rect 338028 5510 338080 5516
rect 335372 3454 336320 3482
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3454
rect 337476 3324 337528 3330
rect 337476 3266 337528 3272
rect 337488 480 337516 3266
rect 338684 480 338712 8978
rect 339328 5642 339356 57530
rect 339420 5710 339448 59758
rect 340156 59758 340194 59786
rect 341066 59786 341094 60044
rect 341966 59786 341994 60044
rect 342886 59786 342914 60044
rect 343786 59786 343814 60044
rect 344686 59786 344714 60044
rect 345586 59786 345614 60044
rect 341066 59758 341104 59786
rect 341966 59758 342208 59786
rect 342886 59758 342944 59786
rect 343786 59758 343864 59786
rect 344686 59758 344876 59786
rect 340052 57792 340104 57798
rect 340052 57734 340104 57740
rect 340064 55214 340092 57734
rect 340156 57594 340184 59758
rect 341076 57594 341104 59758
rect 340144 57588 340196 57594
rect 340144 57530 340196 57536
rect 340788 57588 340840 57594
rect 340788 57530 340840 57536
rect 341064 57588 341116 57594
rect 341064 57530 341116 57536
rect 342076 57588 342128 57594
rect 342076 57530 342128 57536
rect 340064 55186 340184 55214
rect 340156 9042 340184 55186
rect 340144 9036 340196 9042
rect 340144 8978 340196 8984
rect 340800 6594 340828 57530
rect 340880 12232 340932 12238
rect 340880 12174 340932 12180
rect 340788 6588 340840 6594
rect 340788 6530 340840 6536
rect 339408 5704 339460 5710
rect 339408 5646 339460 5652
rect 339316 5636 339368 5642
rect 339316 5578 339368 5584
rect 339868 5568 339920 5574
rect 339868 5510 339920 5516
rect 339880 480 339908 5510
rect 340892 1970 340920 12174
rect 342088 6118 342116 57530
rect 342076 6112 342128 6118
rect 342076 6054 342128 6060
rect 342180 5778 342208 59758
rect 342916 57594 342944 59758
rect 343836 57730 343864 59758
rect 343824 57724 343876 57730
rect 343824 57666 343876 57672
rect 342904 57588 342956 57594
rect 342904 57530 342956 57536
rect 343548 57588 343600 57594
rect 343548 57530 343600 57536
rect 342904 57180 342956 57186
rect 342904 57122 342956 57128
rect 342168 5772 342220 5778
rect 342168 5714 342220 5720
rect 340972 4072 341024 4078
rect 340972 4014 341024 4020
rect 340880 1964 340932 1970
rect 340880 1906 340932 1912
rect 340984 480 341012 4014
rect 342916 3874 342944 57122
rect 343560 5846 343588 57530
rect 344848 5982 344876 59758
rect 345584 59758 345614 59786
rect 346486 59786 346514 60044
rect 347386 59786 347414 60044
rect 348286 59786 348314 60044
rect 349206 59786 349234 60044
rect 350106 59786 350134 60044
rect 351006 59786 351034 60044
rect 351906 59786 351934 60044
rect 352806 59786 352834 60044
rect 353706 59786 353734 60044
rect 354606 59786 354634 60044
rect 355526 59786 355554 60044
rect 346486 59758 346532 59786
rect 347386 59758 347636 59786
rect 348286 59758 348372 59786
rect 349206 59758 349292 59786
rect 350106 59758 350488 59786
rect 351006 59758 351040 59786
rect 351906 59758 351960 59786
rect 352806 59758 353156 59786
rect 345584 57730 345612 59758
rect 346504 57730 346532 59758
rect 344928 57724 344980 57730
rect 344928 57666 344980 57672
rect 345572 57724 345624 57730
rect 345572 57666 345624 57672
rect 346308 57724 346360 57730
rect 346308 57666 346360 57672
rect 346492 57724 346544 57730
rect 346492 57666 346544 57672
rect 344836 5976 344888 5982
rect 344836 5918 344888 5924
rect 344940 5914 344968 57666
rect 345664 56296 345716 56302
rect 345664 56238 345716 56244
rect 345020 21480 345072 21486
rect 345020 21422 345072 21428
rect 345032 16574 345060 21422
rect 345032 16546 345336 16574
rect 344928 5908 344980 5914
rect 344928 5850 344980 5856
rect 343548 5840 343600 5846
rect 343548 5782 343600 5788
rect 343364 5636 343416 5642
rect 343364 5578 343416 5584
rect 342904 3868 342956 3874
rect 342904 3810 342956 3816
rect 342168 1964 342220 1970
rect 342168 1906 342220 1912
rect 342180 480 342208 1906
rect 343376 480 343404 5578
rect 344560 4140 344612 4146
rect 344560 4082 344612 4088
rect 344572 480 344600 4082
rect 345308 490 345336 16546
rect 345676 3330 345704 56238
rect 346320 6050 346348 57666
rect 347608 6866 347636 59758
rect 348344 57730 348372 59758
rect 349264 57730 349292 59758
rect 347688 57724 347740 57730
rect 347688 57666 347740 57672
rect 348332 57724 348384 57730
rect 348332 57666 348384 57672
rect 349068 57724 349120 57730
rect 349068 57666 349120 57672
rect 349252 57724 349304 57730
rect 349252 57666 349304 57672
rect 350356 57724 350408 57730
rect 350356 57666 350408 57672
rect 347596 6860 347648 6866
rect 347596 6802 347648 6808
rect 347700 6118 347728 57666
rect 349080 6798 349108 57666
rect 349252 13524 349304 13530
rect 349252 13466 349304 13472
rect 349068 6792 349120 6798
rect 349068 6734 349120 6740
rect 347688 6112 347740 6118
rect 347688 6054 347740 6060
rect 346308 6044 346360 6050
rect 346308 5986 346360 5992
rect 346952 5704 347004 5710
rect 346952 5646 347004 5652
rect 345664 3324 345716 3330
rect 345664 3266 345716 3272
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 5646
rect 348056 3324 348108 3330
rect 348056 3266 348108 3272
rect 348068 480 348096 3266
rect 349264 480 349292 13466
rect 350368 6730 350396 57666
rect 350356 6724 350408 6730
rect 350356 6666 350408 6672
rect 350460 6662 350488 59758
rect 351012 57730 351040 59758
rect 351932 57730 351960 59758
rect 351000 57724 351052 57730
rect 351000 57666 351052 57672
rect 351828 57724 351880 57730
rect 351828 57666 351880 57672
rect 351920 57724 351972 57730
rect 351920 57666 351972 57672
rect 350448 6656 350500 6662
rect 350448 6598 350500 6604
rect 351840 6594 351868 57666
rect 352840 9036 352892 9042
rect 352840 8978 352892 8984
rect 350356 6588 350408 6594
rect 350356 6530 350408 6536
rect 351828 6588 351880 6594
rect 351828 6530 351880 6536
rect 350368 626 350396 6530
rect 351642 3360 351698 3369
rect 351642 3295 351698 3304
rect 350368 598 350488 626
rect 350460 480 350488 598
rect 351656 480 351684 3295
rect 352852 480 352880 8978
rect 353128 7070 353156 59758
rect 353680 59758 353734 59786
rect 354600 59758 354634 59786
rect 355520 59758 355554 59786
rect 356426 59786 356454 60044
rect 357326 59786 357354 60044
rect 358226 59786 358254 60044
rect 359126 59786 359154 60044
rect 356426 59758 356468 59786
rect 357326 59758 357388 59786
rect 358226 59758 358308 59786
rect 353680 57866 353708 59758
rect 353668 57860 353720 57866
rect 353668 57802 353720 57808
rect 353208 57724 353260 57730
rect 353208 57666 353260 57672
rect 353944 57724 353996 57730
rect 353944 57666 353996 57672
rect 353116 7064 353168 7070
rect 353116 7006 353168 7012
rect 353220 5574 353248 57666
rect 353956 16574 353984 57666
rect 353864 16546 353984 16574
rect 353864 8974 353892 16546
rect 353944 13524 353996 13530
rect 353944 13466 353996 13472
rect 353852 8968 353904 8974
rect 353852 8910 353904 8916
rect 353208 5568 353260 5574
rect 353208 5510 353260 5516
rect 353956 3398 353984 13466
rect 354600 12306 354628 59758
rect 355520 57934 355548 59758
rect 355508 57928 355560 57934
rect 355508 57870 355560 57876
rect 356440 57798 356468 59758
rect 356428 57792 356480 57798
rect 356428 57734 356480 57740
rect 357256 57792 357308 57798
rect 357256 57734 357308 57740
rect 356336 13388 356388 13394
rect 356336 13330 356388 13336
rect 354588 12300 354640 12306
rect 354588 12242 354640 12248
rect 354036 5704 354088 5710
rect 354036 5646 354088 5652
rect 353944 3392 353996 3398
rect 353944 3334 353996 3340
rect 354048 480 354076 5646
rect 355230 3496 355286 3505
rect 355230 3431 355286 3440
rect 355244 480 355272 3431
rect 356348 480 356376 13330
rect 357268 8430 357296 57734
rect 357360 8498 357388 59758
rect 358084 57928 358136 57934
rect 358084 57870 358136 57876
rect 358096 17542 358124 57870
rect 358280 57798 358308 59758
rect 359108 59758 359154 59786
rect 360026 59786 360054 60044
rect 360946 59786 360974 60044
rect 361846 59786 361874 60044
rect 362746 59786 362774 60044
rect 363646 59786 363674 60044
rect 364546 59786 364574 60044
rect 360026 59758 360056 59786
rect 360946 59758 360976 59786
rect 361846 59758 361896 59786
rect 362746 59758 362816 59786
rect 359108 57798 359136 59758
rect 358268 57792 358320 57798
rect 358268 57734 358320 57740
rect 358728 57792 358780 57798
rect 358728 57734 358780 57740
rect 359096 57792 359148 57798
rect 359096 57734 359148 57740
rect 358084 17536 358136 17542
rect 358084 17478 358136 17484
rect 358176 17468 358228 17474
rect 358176 17410 358228 17416
rect 357348 8492 357400 8498
rect 357348 8434 357400 8440
rect 357256 8424 357308 8430
rect 357256 8366 357308 8372
rect 357532 5772 357584 5778
rect 357532 5714 357584 5720
rect 357544 480 357572 5714
rect 358188 3806 358216 17410
rect 358740 8566 358768 57734
rect 359464 12096 359516 12102
rect 359464 12038 359516 12044
rect 358728 8560 358780 8566
rect 358728 8502 358780 8508
rect 358176 3800 358228 3806
rect 358176 3742 358228 3748
rect 358726 3632 358782 3641
rect 358726 3567 358782 3576
rect 358740 480 358768 3567
rect 359476 490 359504 12038
rect 360028 8702 360056 59758
rect 360948 57798 360976 59758
rect 361868 57798 361896 59758
rect 360108 57792 360160 57798
rect 360108 57734 360160 57740
rect 360936 57792 360988 57798
rect 360936 57734 360988 57740
rect 361488 57792 361540 57798
rect 361488 57734 361540 57740
rect 361856 57792 361908 57798
rect 361856 57734 361908 57740
rect 360016 8696 360068 8702
rect 360016 8638 360068 8644
rect 360120 8634 360148 57734
rect 360844 32428 360896 32434
rect 360844 32370 360896 32376
rect 360108 8628 360160 8634
rect 360108 8570 360160 8576
rect 360856 3942 360884 32370
rect 361500 8770 361528 57734
rect 362788 8906 362816 59758
rect 363616 59758 363674 59786
rect 364536 59758 364574 59786
rect 365446 59786 365474 60044
rect 366346 59786 366374 60044
rect 367266 59786 367294 60044
rect 368166 59786 368194 60044
rect 369066 59786 369094 60044
rect 369966 59786 369994 60044
rect 365446 59758 365668 59786
rect 366346 59758 366404 59786
rect 367266 59758 367324 59786
rect 368166 59758 368336 59786
rect 363616 57934 363644 59758
rect 363604 57928 363656 57934
rect 363604 57870 363656 57876
rect 364248 57928 364300 57934
rect 364248 57870 364300 57876
rect 362868 57792 362920 57798
rect 362868 57734 362920 57740
rect 363604 57792 363656 57798
rect 363604 57734 363656 57740
rect 362776 8900 362828 8906
rect 362776 8842 362828 8848
rect 362880 8838 362908 57734
rect 362868 8832 362920 8838
rect 362868 8774 362920 8780
rect 361488 8764 361540 8770
rect 361488 8706 361540 8712
rect 363512 6520 363564 6526
rect 363512 6462 363564 6468
rect 361120 5840 361172 5846
rect 361120 5782 361172 5788
rect 360844 3936 360896 3942
rect 360844 3878 360896 3884
rect 359752 598 359964 626
rect 359752 490 359780 598
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 462 359780 490
rect 359936 480 359964 598
rect 361132 480 361160 5782
rect 362314 3768 362370 3777
rect 362314 3703 362370 3712
rect 362328 480 362356 3703
rect 363524 480 363552 6462
rect 363616 4010 363644 57734
rect 364260 9654 364288 57870
rect 364536 57662 364564 59758
rect 364524 57656 364576 57662
rect 364524 57598 364576 57604
rect 365536 57656 365588 57662
rect 365536 57598 365588 57604
rect 364248 9648 364300 9654
rect 364248 9590 364300 9596
rect 365548 9586 365576 57598
rect 365536 9580 365588 9586
rect 365536 9522 365588 9528
rect 365640 9518 365668 59758
rect 366376 57662 366404 59758
rect 367296 57662 367324 59758
rect 366364 57656 366416 57662
rect 366364 57598 366416 57604
rect 367008 57656 367060 57662
rect 367008 57598 367060 57604
rect 367284 57656 367336 57662
rect 367284 57598 367336 57604
rect 365628 9512 365680 9518
rect 365628 9454 365680 9460
rect 367020 9450 367048 57598
rect 367008 9444 367060 9450
rect 367008 9386 367060 9392
rect 368308 9314 368336 59758
rect 369044 59758 369094 59786
rect 369964 59758 369994 59786
rect 370866 59786 370894 60044
rect 371766 59786 371794 60044
rect 372666 59786 372694 60044
rect 373586 59786 373614 60044
rect 374486 59786 374514 60044
rect 370866 59758 371096 59786
rect 371766 59758 371832 59786
rect 372666 59758 372752 59786
rect 373586 59758 373672 59786
rect 369044 57662 369072 59758
rect 369964 57662 369992 59758
rect 368388 57656 368440 57662
rect 368388 57598 368440 57604
rect 369032 57656 369084 57662
rect 369032 57598 369084 57604
rect 369768 57656 369820 57662
rect 369768 57598 369820 57604
rect 369952 57656 370004 57662
rect 369952 57598 370004 57604
rect 368400 9382 368428 57598
rect 368388 9376 368440 9382
rect 368388 9318 368440 9324
rect 368296 9308 368348 9314
rect 368296 9250 368348 9256
rect 369780 9246 369808 57598
rect 369768 9240 369820 9246
rect 369768 9182 369820 9188
rect 371068 9110 371096 59758
rect 371804 57662 371832 59758
rect 372724 57662 372752 59758
rect 371148 57656 371200 57662
rect 371148 57598 371200 57604
rect 371792 57656 371844 57662
rect 371792 57598 371844 57604
rect 372528 57656 372580 57662
rect 372528 57598 372580 57604
rect 372712 57656 372764 57662
rect 372712 57598 372764 57604
rect 371160 9178 371188 57598
rect 371884 57180 371936 57186
rect 371884 57122 371936 57128
rect 371148 9172 371200 9178
rect 371148 9114 371200 9120
rect 371056 9104 371108 9110
rect 371056 9046 371108 9052
rect 367008 6452 367060 6458
rect 367008 6394 367060 6400
rect 364616 5908 364668 5914
rect 364616 5850 364668 5856
rect 363604 4004 363656 4010
rect 363604 3946 363656 3952
rect 364628 480 364656 5850
rect 365812 3800 365864 3806
rect 365812 3742 365864 3748
rect 365824 480 365852 3742
rect 367020 480 367048 6394
rect 371896 6390 371924 57122
rect 372540 9042 372568 57598
rect 373644 56710 373672 59758
rect 374472 59758 374514 59786
rect 375386 59786 375414 60044
rect 376286 59786 376314 60044
rect 377186 59786 377214 60044
rect 378086 59786 378114 60044
rect 379006 59786 379034 60044
rect 379906 59786 379934 60044
rect 375386 59758 375420 59786
rect 376286 59758 376708 59786
rect 377186 59758 377260 59786
rect 374472 57662 374500 59758
rect 375392 57662 375420 59758
rect 373908 57656 373960 57662
rect 373908 57598 373960 57604
rect 374460 57656 374512 57662
rect 374460 57598 374512 57604
rect 375288 57656 375340 57662
rect 375288 57598 375340 57604
rect 375380 57656 375432 57662
rect 375380 57598 375432 57604
rect 376576 57656 376628 57662
rect 376576 57598 376628 57604
rect 373632 56704 373684 56710
rect 373632 56646 373684 56652
rect 372528 9036 372580 9042
rect 372528 8978 372580 8984
rect 373920 8974 373948 57598
rect 374644 56704 374696 56710
rect 374644 56646 374696 56652
rect 374656 29646 374684 56646
rect 374644 29640 374696 29646
rect 374644 29582 374696 29588
rect 374644 20052 374696 20058
rect 374644 19994 374696 20000
rect 373908 8968 373960 8974
rect 373908 8910 373960 8916
rect 370596 6384 370648 6390
rect 370596 6326 370648 6332
rect 371884 6384 371936 6390
rect 371884 6326 371936 6332
rect 368204 5976 368256 5982
rect 368204 5918 368256 5924
rect 368216 480 368244 5918
rect 369400 3868 369452 3874
rect 369400 3810 369452 3816
rect 369412 480 369440 3810
rect 370608 480 370636 6326
rect 374092 6316 374144 6322
rect 374092 6258 374144 6264
rect 371700 6044 371752 6050
rect 371700 5986 371752 5992
rect 371712 480 371740 5986
rect 372896 3936 372948 3942
rect 372896 3878 372948 3884
rect 372908 480 372936 3878
rect 374104 480 374132 6258
rect 374656 3330 374684 19994
rect 375300 12238 375328 57598
rect 376588 25566 376616 57598
rect 376576 25560 376628 25566
rect 376576 25502 376628 25508
rect 376024 22840 376076 22846
rect 376024 22782 376076 22788
rect 375288 12232 375340 12238
rect 375288 12174 375340 12180
rect 375288 6112 375340 6118
rect 375288 6054 375340 6060
rect 374644 3324 374696 3330
rect 374644 3266 374696 3272
rect 375300 480 375328 6054
rect 376036 4078 376064 22782
rect 376680 12102 376708 59758
rect 377232 57662 377260 59758
rect 378060 59758 378114 59786
rect 378980 59758 379034 59786
rect 379900 59758 379934 59786
rect 380806 59786 380834 60044
rect 381706 59786 381734 60044
rect 382606 59786 382634 60044
rect 383506 59786 383534 60044
rect 384406 59786 384434 60044
rect 385326 59786 385354 60044
rect 386226 59786 386254 60044
rect 387126 59786 387154 60044
rect 388026 59786 388054 60044
rect 380806 59758 380848 59786
rect 381706 59758 381768 59786
rect 382606 59758 382688 59786
rect 383506 59758 383608 59786
rect 384406 59758 384436 59786
rect 385326 59758 385356 59786
rect 386226 59758 386276 59786
rect 387126 59758 387196 59786
rect 377220 57656 377272 57662
rect 377220 57598 377272 57604
rect 377956 57656 378008 57662
rect 377956 57598 378008 57604
rect 377968 16250 377996 57598
rect 377956 16244 378008 16250
rect 377956 16186 378008 16192
rect 377404 14884 377456 14890
rect 377404 14826 377456 14832
rect 376668 12096 376720 12102
rect 376668 12038 376720 12044
rect 377416 4146 377444 14826
rect 378060 13394 378088 59758
rect 378784 57860 378836 57866
rect 378784 57802 378836 57808
rect 378048 13388 378100 13394
rect 378048 13330 378100 13336
rect 378796 12374 378824 57802
rect 378980 57662 379008 59758
rect 379900 57934 379928 59758
rect 379888 57928 379940 57934
rect 379888 57870 379940 57876
rect 378968 57656 379020 57662
rect 378968 57598 379020 57604
rect 379428 57656 379480 57662
rect 379428 57598 379480 57604
rect 379440 13598 379468 57598
rect 380820 56234 380848 59758
rect 381544 57860 381596 57866
rect 381544 57802 381596 57808
rect 380808 56228 380860 56234
rect 380808 56170 380860 56176
rect 379428 13592 379480 13598
rect 379428 13534 379480 13540
rect 378784 12368 378836 12374
rect 378784 12310 378836 12316
rect 381556 11762 381584 57802
rect 381740 57662 381768 59758
rect 382660 57662 382688 59758
rect 381728 57656 381780 57662
rect 381728 57598 381780 57604
rect 382188 57656 382240 57662
rect 382188 57598 382240 57604
rect 382648 57656 382700 57662
rect 382648 57598 382700 57604
rect 383476 57656 383528 57662
rect 383476 57598 383528 57604
rect 381544 11756 381596 11762
rect 381544 11698 381596 11704
rect 378876 6860 378928 6866
rect 378876 6802 378928 6808
rect 377680 6248 377732 6254
rect 377680 6190 377732 6196
rect 377404 4140 377456 4146
rect 377404 4082 377456 4088
rect 376024 4072 376076 4078
rect 376024 4014 376076 4020
rect 376484 4004 376536 4010
rect 376484 3946 376536 3952
rect 376496 480 376524 3946
rect 377692 480 377720 6190
rect 378888 480 378916 6802
rect 381176 6180 381228 6186
rect 381176 6122 381228 6128
rect 379980 4072 380032 4078
rect 379980 4014 380032 4020
rect 379992 480 380020 4014
rect 381188 480 381216 6122
rect 382200 5642 382228 57598
rect 382372 6792 382424 6798
rect 382372 6734 382424 6740
rect 382188 5636 382240 5642
rect 382188 5578 382240 5584
rect 382384 480 382412 6734
rect 383488 5710 383516 57598
rect 383580 5778 383608 59758
rect 384408 57526 384436 59758
rect 385328 57526 385356 59758
rect 384396 57520 384448 57526
rect 384396 57462 384448 57468
rect 384948 57520 385000 57526
rect 384948 57462 385000 57468
rect 385316 57520 385368 57526
rect 385316 57462 385368 57468
rect 384764 6384 384816 6390
rect 384764 6326 384816 6332
rect 383568 5772 383620 5778
rect 383568 5714 383620 5720
rect 383476 5704 383528 5710
rect 383476 5646 383528 5652
rect 383568 4140 383620 4146
rect 383568 4082 383620 4088
rect 383580 480 383608 4082
rect 384776 480 384804 6326
rect 384960 6050 384988 57462
rect 385960 6724 386012 6730
rect 385960 6666 386012 6672
rect 384948 6044 385000 6050
rect 384948 5986 385000 5992
rect 385972 480 386000 6666
rect 386248 5982 386276 59758
rect 387168 57526 387196 59758
rect 387996 59758 388054 59786
rect 388926 59786 388954 60044
rect 389826 59786 389854 60044
rect 390726 59786 390754 60044
rect 391646 59786 391674 60044
rect 392546 59786 392574 60044
rect 393446 59786 393474 60044
rect 388926 59758 389036 59786
rect 389826 59758 389864 59786
rect 390726 59758 390784 59786
rect 391646 59758 391796 59786
rect 392546 59758 392624 59786
rect 387996 57526 388024 59758
rect 386328 57520 386380 57526
rect 386328 57462 386380 57468
rect 387156 57520 387208 57526
rect 387156 57462 387208 57468
rect 387708 57520 387760 57526
rect 387708 57462 387760 57468
rect 387984 57520 388036 57526
rect 387984 57462 388036 57468
rect 386236 5976 386288 5982
rect 386236 5918 386288 5924
rect 386340 5914 386368 57462
rect 387720 6186 387748 57462
rect 387800 13252 387852 13258
rect 387800 13194 387852 13200
rect 387708 6180 387760 6186
rect 387708 6122 387760 6128
rect 386328 5908 386380 5914
rect 386328 5850 386380 5856
rect 387156 3392 387208 3398
rect 387156 3334 387208 3340
rect 387168 480 387196 3334
rect 387812 490 387840 13194
rect 389008 6254 389036 59758
rect 389836 57526 389864 59758
rect 390756 57526 390784 59758
rect 389088 57520 389140 57526
rect 389088 57462 389140 57468
rect 389824 57520 389876 57526
rect 389824 57462 389876 57468
rect 390468 57520 390520 57526
rect 390468 57462 390520 57468
rect 390744 57520 390796 57526
rect 390744 57462 390796 57468
rect 388996 6248 389048 6254
rect 388996 6190 389048 6196
rect 389100 6118 389128 57462
rect 389824 57180 389876 57186
rect 389824 57122 389876 57128
rect 389836 6866 389864 57122
rect 389824 6860 389876 6866
rect 389824 6802 389876 6808
rect 390480 6798 390508 57462
rect 391768 12434 391796 59758
rect 392596 57526 392624 59758
rect 393424 59758 393474 59786
rect 394346 59786 394374 60044
rect 395246 59786 395274 60044
rect 396146 59786 396174 60044
rect 397066 59786 397094 60044
rect 397966 59786 397994 60044
rect 398866 59786 398894 60044
rect 399766 59786 399794 60044
rect 394346 59758 394556 59786
rect 395246 59758 395292 59786
rect 396146 59758 396212 59786
rect 397066 59758 397408 59786
rect 397966 59758 398052 59786
rect 398866 59758 398972 59786
rect 392676 57928 392728 57934
rect 392676 57870 392728 57876
rect 391848 57520 391900 57526
rect 391848 57462 391900 57468
rect 392584 57520 392636 57526
rect 392584 57462 392636 57468
rect 391676 12406 391796 12434
rect 390468 6792 390520 6798
rect 390468 6734 390520 6740
rect 391676 6662 391704 12406
rect 391860 9602 391888 57462
rect 392688 45554 392716 57870
rect 393424 57526 393452 59758
rect 393228 57520 393280 57526
rect 393228 57462 393280 57468
rect 393412 57520 393464 57526
rect 393412 57462 393464 57468
rect 392596 45526 392716 45554
rect 392596 17270 392624 45526
rect 392584 17264 392636 17270
rect 392584 17206 392636 17212
rect 391768 9574 391888 9602
rect 391768 6730 391796 9574
rect 391848 6860 391900 6866
rect 391848 6802 391900 6808
rect 391756 6724 391808 6730
rect 391756 6666 391808 6672
rect 389456 6656 389508 6662
rect 389456 6598 389508 6604
rect 391664 6656 391716 6662
rect 391664 6598 391716 6604
rect 389088 6112 389140 6118
rect 389088 6054 389140 6060
rect 388088 598 388300 626
rect 388088 490 388116 598
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 462 388116 490
rect 388272 480 388300 598
rect 389468 480 389496 6598
rect 390652 3324 390704 3330
rect 390652 3266 390704 3272
rect 390664 480 390692 3266
rect 391860 480 391888 6802
rect 393240 6594 393268 57462
rect 393044 6588 393096 6594
rect 393044 6530 393096 6536
rect 393228 6588 393280 6594
rect 393228 6530 393280 6536
rect 393056 480 393084 6530
rect 394528 6458 394556 59758
rect 395264 57526 395292 59758
rect 396184 57526 396212 59758
rect 394608 57520 394660 57526
rect 394608 57462 394660 57468
rect 395252 57520 395304 57526
rect 395252 57462 395304 57468
rect 395988 57520 396040 57526
rect 395988 57462 396040 57468
rect 396172 57520 396224 57526
rect 396172 57462 396224 57468
rect 397276 57520 397328 57526
rect 397276 57462 397328 57468
rect 394620 6526 394648 57462
rect 394700 22772 394752 22778
rect 394700 22714 394752 22720
rect 394712 16574 394740 22714
rect 394712 16546 395384 16574
rect 394608 6520 394660 6526
rect 394608 6462 394660 6468
rect 394516 6452 394568 6458
rect 394516 6394 394568 6400
rect 394240 3256 394292 3262
rect 394240 3198 394292 3204
rect 394252 480 394280 3198
rect 395356 480 395384 16546
rect 396000 6390 396028 57462
rect 395988 6384 396040 6390
rect 395988 6326 396040 6332
rect 397288 6322 397316 57462
rect 396540 6316 396592 6322
rect 396540 6258 396592 6264
rect 397276 6316 397328 6322
rect 397276 6258 397328 6264
rect 396552 480 396580 6258
rect 397380 6254 397408 59758
rect 398024 57526 398052 59758
rect 398012 57520 398064 57526
rect 398012 57462 398064 57468
rect 398748 57520 398800 57526
rect 398748 57462 398800 57468
rect 397368 6248 397420 6254
rect 397368 6190 397420 6196
rect 398760 6186 398788 57462
rect 398840 14680 398892 14686
rect 398840 14622 398892 14628
rect 398852 6914 398880 14622
rect 398944 10334 398972 59758
rect 399036 59758 399794 59786
rect 400666 59786 400694 60044
rect 401566 59786 401594 60044
rect 402466 59786 402494 60044
rect 400666 59758 400720 59786
rect 401566 59758 401640 59786
rect 399036 10402 399064 59758
rect 400692 57866 400720 59758
rect 400680 57860 400732 57866
rect 400680 57802 400732 57808
rect 401612 57526 401640 59758
rect 402440 59758 402494 59786
rect 402980 59832 403032 59838
rect 403386 59786 403414 60044
rect 404286 59838 404314 60044
rect 402980 59774 403032 59780
rect 402440 57934 402468 59758
rect 402428 57928 402480 57934
rect 402428 57870 402480 57876
rect 400864 57520 400916 57526
rect 400864 57462 400916 57468
rect 401600 57520 401652 57526
rect 401600 57462 401652 57468
rect 401692 57520 401744 57526
rect 401692 57462 401744 57468
rect 400876 15910 400904 57462
rect 401704 57338 401732 57462
rect 401520 57310 401732 57338
rect 400864 15904 400916 15910
rect 400864 15846 400916 15852
rect 399024 10396 399076 10402
rect 399024 10338 399076 10344
rect 398932 10328 398984 10334
rect 398932 10270 398984 10276
rect 400128 7064 400180 7070
rect 400128 7006 400180 7012
rect 398852 6886 398972 6914
rect 398748 6180 398800 6186
rect 398748 6122 398800 6128
rect 397736 3188 397788 3194
rect 397736 3130 397788 3136
rect 397748 480 397776 3130
rect 398944 480 398972 6886
rect 400140 480 400168 7006
rect 401520 6914 401548 57310
rect 402520 11960 402572 11966
rect 402520 11902 402572 11908
rect 401336 6886 401548 6914
rect 401336 480 401364 6886
rect 402532 480 402560 11902
rect 402992 3534 403020 59774
rect 403084 59758 403414 59786
rect 404274 59832 404326 59838
rect 405186 59786 405214 60044
rect 404274 59774 404326 59780
rect 404372 59758 405214 59786
rect 405740 59832 405792 59838
rect 406086 59786 406114 60044
rect 406986 59838 407014 60044
rect 405740 59774 405792 59780
rect 402980 3528 403032 3534
rect 402980 3470 403032 3476
rect 403084 3466 403112 59758
rect 403624 12368 403676 12374
rect 403624 12310 403676 12316
rect 403072 3460 403124 3466
rect 403072 3402 403124 3408
rect 403636 480 403664 12310
rect 404372 3602 404400 59758
rect 405752 3738 405780 59774
rect 405844 59758 406114 59786
rect 406974 59832 407026 59838
rect 407886 59786 407914 60044
rect 408786 59786 408814 60044
rect 409706 59786 409734 60044
rect 410606 59786 410634 60044
rect 406974 59774 407026 59780
rect 407224 59758 407914 59786
rect 408512 59758 408814 59786
rect 408972 59758 409734 59786
rect 409892 59758 410634 59786
rect 411260 59832 411312 59838
rect 411506 59786 411534 60044
rect 412406 59838 412434 60044
rect 411260 59774 411312 59780
rect 405740 3732 405792 3738
rect 405740 3674 405792 3680
rect 405844 3670 405872 59758
rect 406016 14612 406068 14618
rect 406016 14554 406068 14560
rect 405832 3664 405884 3670
rect 405832 3606 405884 3612
rect 404360 3596 404412 3602
rect 404360 3538 404412 3544
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 404832 480 404860 3402
rect 406028 480 406056 14554
rect 407120 12300 407172 12306
rect 407120 12242 407172 12248
rect 407132 6914 407160 12242
rect 407224 10470 407252 59758
rect 407764 57452 407816 57458
rect 407764 57394 407816 57400
rect 407212 10464 407264 10470
rect 407212 10406 407264 10412
rect 407132 6886 407252 6914
rect 407224 480 407252 6886
rect 407776 4214 407804 57394
rect 408512 10538 408540 59758
rect 408972 45554 409000 59758
rect 408604 45526 409000 45554
rect 408604 10606 408632 45526
rect 409892 10674 409920 59758
rect 410524 57452 410576 57458
rect 410524 57394 410576 57400
rect 410536 19990 410564 57394
rect 410524 19984 410576 19990
rect 410524 19926 410576 19932
rect 409972 17536 410024 17542
rect 409972 17478 410024 17484
rect 409984 16574 410012 17478
rect 409984 16546 410840 16574
rect 409880 10668 409932 10674
rect 409880 10610 409932 10616
rect 408592 10600 408644 10606
rect 408592 10542 408644 10548
rect 408500 10532 408552 10538
rect 408500 10474 408552 10480
rect 407764 4208 407816 4214
rect 407764 4150 407816 4156
rect 409604 4208 409656 4214
rect 409604 4150 409656 4156
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 409616 480 409644 4150
rect 410812 480 410840 16546
rect 411272 10810 411300 59774
rect 411364 59758 411534 59786
rect 412394 59832 412446 59838
rect 413306 59786 413334 60044
rect 412394 59774 412446 59780
rect 412652 59758 413334 59786
rect 414020 59832 414072 59838
rect 414206 59786 414234 60044
rect 415126 59838 415154 60044
rect 414020 59774 414072 59780
rect 411260 10804 411312 10810
rect 411260 10746 411312 10752
rect 411364 10742 411392 59758
rect 412652 10878 412680 59758
rect 412732 24132 412784 24138
rect 412732 24074 412784 24080
rect 412640 10872 412692 10878
rect 412640 10814 412692 10820
rect 411352 10736 411404 10742
rect 411352 10678 411404 10684
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 412744 490 412772 24074
rect 414032 11014 414060 59774
rect 414124 59758 414234 59786
rect 415114 59832 415166 59838
rect 416026 59786 416054 60044
rect 415114 59774 415166 59780
rect 415412 59758 416054 59786
rect 416780 59832 416832 59838
rect 416926 59786 416954 60044
rect 417826 59838 417854 60044
rect 416780 59774 416832 59780
rect 414020 11008 414072 11014
rect 414020 10950 414072 10956
rect 414124 10946 414152 59758
rect 414112 10940 414164 10946
rect 414112 10882 414164 10888
rect 415412 10266 415440 59758
rect 415400 10260 415452 10266
rect 415400 10202 415452 10208
rect 416792 10130 416820 59774
rect 416884 59758 416954 59786
rect 417814 59832 417866 59838
rect 418726 59786 418754 60044
rect 417814 59774 417866 59780
rect 418172 59758 418754 59786
rect 419540 59832 419592 59838
rect 419540 59774 419592 59780
rect 419626 59786 419654 60044
rect 420526 59838 420554 60044
rect 420514 59832 420566 59838
rect 416884 10198 416912 59758
rect 416872 10192 416924 10198
rect 416872 10134 416924 10140
rect 416780 10124 416832 10130
rect 416780 10066 416832 10072
rect 418172 10062 418200 59758
rect 418804 57656 418856 57662
rect 418804 57598 418856 57604
rect 418816 10334 418844 57598
rect 418804 10328 418856 10334
rect 418804 10270 418856 10276
rect 418160 10056 418212 10062
rect 418160 9998 418212 10004
rect 419552 9926 419580 59774
rect 419626 59758 419672 59786
rect 421446 59786 421474 60044
rect 422346 59786 422374 60044
rect 423246 59786 423274 60044
rect 424146 59786 424174 60044
rect 420514 59774 420566 59780
rect 419644 9994 419672 59758
rect 420932 59758 421474 59786
rect 422312 59758 422374 59786
rect 423232 59758 423274 59786
rect 423692 59758 424174 59786
rect 425046 59786 425074 60044
rect 425946 59786 425974 60044
rect 426846 59786 426874 60044
rect 427766 59786 427794 60044
rect 428666 59786 428694 60044
rect 425046 59758 425192 59786
rect 420932 15978 420960 59758
rect 422312 56642 422340 59758
rect 423232 57458 423260 59758
rect 423220 57452 423272 57458
rect 423220 57394 423272 57400
rect 423588 57452 423640 57458
rect 423588 57394 423640 57400
rect 421564 56636 421616 56642
rect 421564 56578 421616 56584
rect 422300 56636 422352 56642
rect 422300 56578 422352 56584
rect 421576 18630 421604 56578
rect 421564 18624 421616 18630
rect 421564 18566 421616 18572
rect 420920 15972 420972 15978
rect 420920 15914 420972 15920
rect 419632 9988 419684 9994
rect 419632 9930 419684 9936
rect 419540 9920 419592 9926
rect 419540 9862 419592 9868
rect 421380 8560 421432 8566
rect 421380 8502 421432 8508
rect 417884 8492 417936 8498
rect 417884 8434 417936 8440
rect 414296 8424 414348 8430
rect 414296 8366 414348 8372
rect 412928 598 413140 626
rect 412928 490 412956 598
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412744 462 412956 490
rect 413112 480 413140 598
rect 414308 480 414336 8366
rect 416688 7132 416740 7138
rect 416688 7074 416740 7080
rect 415492 3052 415544 3058
rect 415492 2994 415544 3000
rect 415504 480 415532 2994
rect 416700 480 416728 7074
rect 417896 480 417924 8434
rect 420184 7200 420236 7206
rect 420184 7142 420236 7148
rect 418988 3732 419040 3738
rect 418988 3674 419040 3680
rect 419000 480 419028 3674
rect 420196 480 420224 7142
rect 421392 480 421420 8502
rect 423600 3670 423628 57394
rect 423692 21418 423720 59758
rect 425060 57656 425112 57662
rect 425060 57598 425112 57604
rect 423680 21412 423732 21418
rect 423680 21354 423732 21360
rect 425072 16046 425100 57598
rect 425164 33794 425192 59758
rect 425900 59758 425974 59786
rect 426820 59758 426874 59786
rect 427740 59758 427794 59786
rect 427832 59758 428694 59786
rect 429200 59832 429252 59838
rect 429566 59786 429594 60044
rect 430466 59838 430494 60044
rect 429200 59774 429252 59780
rect 425900 57662 425928 59758
rect 425888 57656 425940 57662
rect 425888 57598 425940 57604
rect 426820 56030 426848 59758
rect 427740 56098 427768 59758
rect 427728 56092 427780 56098
rect 427728 56034 427780 56040
rect 426808 56024 426860 56030
rect 426808 55966 426860 55972
rect 425152 33788 425204 33794
rect 425152 33730 425204 33736
rect 425060 16040 425112 16046
rect 425060 15982 425112 15988
rect 427832 14550 427860 59758
rect 429212 37942 429240 59774
rect 429304 59758 429594 59786
rect 430454 59832 430506 59838
rect 431366 59786 431394 60044
rect 430454 59774 430506 59780
rect 430592 59758 431394 59786
rect 431960 59832 432012 59838
rect 432266 59786 432294 60044
rect 433186 59838 433214 60044
rect 431960 59774 432012 59780
rect 429304 54534 429332 59758
rect 430488 57656 430540 57662
rect 430488 57598 430540 57604
rect 429292 54528 429344 54534
rect 429292 54470 429344 54476
rect 429200 37936 429252 37942
rect 429200 37878 429252 37884
rect 427820 14544 427872 14550
rect 427820 14486 427872 14492
rect 428464 8696 428516 8702
rect 428464 8638 428516 8644
rect 424968 8628 425020 8634
rect 424968 8570 425020 8576
rect 423772 7268 423824 7274
rect 423772 7210 423824 7216
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 423588 3664 423640 3670
rect 423588 3606 423640 3612
rect 422588 480 422616 3606
rect 423784 480 423812 7210
rect 424980 480 425008 8570
rect 427268 7336 427320 7342
rect 427268 7278 427320 7284
rect 426164 3120 426216 3126
rect 426164 3062 426216 3068
rect 426176 480 426204 3062
rect 427280 480 427308 7278
rect 428476 480 428504 8638
rect 430500 3670 430528 57598
rect 430592 17338 430620 59758
rect 431224 57860 431276 57866
rect 431224 57802 431276 57808
rect 430580 17332 430632 17338
rect 430580 17274 430632 17280
rect 431236 13326 431264 57802
rect 431224 13320 431276 13326
rect 431224 13262 431276 13268
rect 431972 13190 432000 59774
rect 432064 59758 432294 59786
rect 433174 59832 433226 59838
rect 433174 59774 433226 59780
rect 434086 59786 434114 60044
rect 434720 59832 434772 59838
rect 434086 59758 434116 59786
rect 434986 59786 435014 60044
rect 435886 59838 435914 60044
rect 434720 59774 434772 59780
rect 432064 36582 432092 59758
rect 434088 56166 434116 59758
rect 434076 56160 434128 56166
rect 434076 56102 434128 56108
rect 432052 36576 432104 36582
rect 432052 36518 432104 36524
rect 434732 14822 434760 59774
rect 434824 59758 435014 59786
rect 435874 59832 435926 59838
rect 436786 59786 436814 60044
rect 437686 59786 437714 60044
rect 435874 59774 435926 59780
rect 436112 59758 436814 59786
rect 437676 59758 437714 59786
rect 438586 59786 438614 60044
rect 439506 59786 439534 60044
rect 438586 59758 438624 59786
rect 434824 28286 434852 59758
rect 434812 28280 434864 28286
rect 434812 28222 434864 28228
rect 436112 16114 436140 59758
rect 437676 57934 437704 59758
rect 437664 57928 437716 57934
rect 437664 57870 437716 57876
rect 438596 57866 438624 59758
rect 438872 59758 439534 59786
rect 440406 59786 440434 60044
rect 441306 59786 441334 60044
rect 442206 59786 442234 60044
rect 440406 59758 440464 59786
rect 436744 57860 436796 57866
rect 436744 57802 436796 57808
rect 438584 57860 438636 57866
rect 438584 57802 438636 57808
rect 436100 16108 436152 16114
rect 436100 16050 436152 16056
rect 434720 14816 434772 14822
rect 434720 14758 434772 14764
rect 431960 13184 432012 13190
rect 431960 13126 432012 13132
rect 436756 12034 436784 57802
rect 438872 17406 438900 59758
rect 440436 57866 440464 59758
rect 440528 59758 441334 59786
rect 441632 59758 442234 59786
rect 443000 59832 443052 59838
rect 443106 59786 443134 60044
rect 444006 59838 444034 60044
rect 443000 59774 443052 59780
rect 439504 57860 439556 57866
rect 439504 57802 439556 57808
rect 440424 57860 440476 57866
rect 440424 57802 440476 57808
rect 438860 17400 438912 17406
rect 438860 17342 438912 17348
rect 439516 14754 439544 57802
rect 440528 54602 440556 59758
rect 441528 57860 441580 57866
rect 441528 57802 441580 57808
rect 440516 54596 440568 54602
rect 440516 54538 440568 54544
rect 439504 14748 439556 14754
rect 439504 14690 439556 14696
rect 436744 12028 436796 12034
rect 436744 11970 436796 11976
rect 439136 8900 439188 8906
rect 439136 8842 439188 8848
rect 435548 8832 435600 8838
rect 435548 8774 435600 8780
rect 432052 8764 432104 8770
rect 432052 8706 432104 8712
rect 430856 7404 430908 7410
rect 430856 7346 430908 7352
rect 429660 3664 429712 3670
rect 429660 3606 429712 3612
rect 430488 3664 430540 3670
rect 430488 3606 430540 3612
rect 429672 480 429700 3606
rect 430868 480 430896 7346
rect 432064 480 432092 8706
rect 434444 7472 434496 7478
rect 434444 7414 434496 7420
rect 433248 2984 433300 2990
rect 433248 2926 433300 2932
rect 433260 480 433288 2926
rect 434456 480 434484 7414
rect 435560 480 435588 8774
rect 437940 7540 437992 7546
rect 437940 7482 437992 7488
rect 436744 2916 436796 2922
rect 436744 2858 436796 2864
rect 436756 480 436784 2858
rect 437952 480 437980 7482
rect 439148 480 439176 8842
rect 441252 8288 441304 8294
rect 441252 8230 441304 8236
rect 440332 2848 440384 2854
rect 440332 2790 440384 2796
rect 440344 480 440372 2790
rect 441264 2774 441292 8230
rect 441540 2854 441568 57802
rect 441632 26926 441660 59758
rect 441620 26920 441672 26926
rect 441620 26862 441672 26868
rect 443012 13462 443040 59774
rect 443104 59758 443134 59786
rect 443994 59832 444046 59838
rect 444906 59786 444934 60044
rect 445826 59922 445854 60044
rect 443994 59774 444046 59780
rect 444852 59758 444934 59786
rect 445772 59894 445854 59922
rect 443104 31074 443132 59758
rect 444852 57594 444880 59758
rect 445772 57730 445800 59894
rect 446726 59786 446754 60044
rect 447626 59786 447654 60044
rect 445864 59758 446754 59786
rect 447152 59758 447654 59786
rect 448526 59786 448554 60044
rect 449426 59786 449454 60044
rect 450326 59786 450354 60044
rect 448526 59758 448652 59786
rect 445760 57724 445812 57730
rect 445760 57666 445812 57672
rect 444840 57588 444892 57594
rect 444840 57530 444892 57536
rect 443092 31068 443144 31074
rect 443092 31010 443144 31016
rect 443000 13456 443052 13462
rect 443000 13398 443052 13404
rect 445864 12170 445892 59758
rect 447152 16182 447180 59758
rect 448520 57588 448572 57594
rect 448520 57530 448572 57536
rect 448428 57384 448480 57390
rect 448428 57326 448480 57332
rect 447140 16176 447192 16182
rect 447140 16118 447192 16124
rect 445852 12164 445904 12170
rect 445852 12106 445904 12112
rect 442632 9648 442684 9654
rect 442632 9590 442684 9596
rect 441528 2848 441580 2854
rect 441528 2790 441580 2796
rect 441264 2746 441476 2774
rect 441448 1442 441476 2746
rect 441448 1414 441568 1442
rect 441540 480 441568 1414
rect 442644 480 442672 9590
rect 446220 9580 446272 9586
rect 446220 9522 446272 9528
rect 445024 8220 445076 8226
rect 445024 8162 445076 8168
rect 443828 2848 443880 2854
rect 443828 2790 443880 2796
rect 443840 480 443868 2790
rect 445036 480 445064 8162
rect 446232 480 446260 9522
rect 448440 2990 448468 57326
rect 448532 13530 448560 57530
rect 448624 17474 448652 59758
rect 449360 59758 449454 59786
rect 449912 59758 450354 59786
rect 451246 59786 451274 60044
rect 452146 59786 452174 60044
rect 451246 59758 451320 59786
rect 449360 57594 449388 59758
rect 449348 57588 449400 57594
rect 449348 57530 449400 57536
rect 449912 32434 449940 59758
rect 451292 57798 451320 59758
rect 452120 59758 452174 59786
rect 452660 59832 452712 59838
rect 453046 59786 453074 60044
rect 453946 59838 453974 60044
rect 452660 59774 452712 59780
rect 451280 57792 451332 57798
rect 451280 57734 451332 57740
rect 450544 57180 450596 57186
rect 450544 57122 450596 57128
rect 449900 32428 449952 32434
rect 449900 32370 449952 32376
rect 448612 17468 448664 17474
rect 448612 17410 448664 17416
rect 448520 13524 448572 13530
rect 448520 13466 448572 13472
rect 449808 9512 449860 9518
rect 449808 9454 449860 9460
rect 448612 8152 448664 8158
rect 448612 8094 448664 8100
rect 447416 2984 447468 2990
rect 447416 2926 447468 2932
rect 448428 2984 448480 2990
rect 448428 2926 448480 2932
rect 447428 480 447456 2926
rect 448624 480 448652 8094
rect 449820 480 449848 9454
rect 450556 8158 450584 57122
rect 452120 56302 452148 59758
rect 452108 56296 452160 56302
rect 452108 56238 452160 56244
rect 452672 14890 452700 59774
rect 452764 59758 453074 59786
rect 453934 59832 453986 59838
rect 454846 59786 454874 60044
rect 455746 59786 455774 60044
rect 456646 59786 456674 60044
rect 457566 59786 457594 60044
rect 458466 59786 458494 60044
rect 459366 59786 459394 60044
rect 460266 59786 460294 60044
rect 461166 59786 461194 60044
rect 462066 59786 462094 60044
rect 462966 59786 462994 60044
rect 453934 59774 453986 59780
rect 454052 59758 454874 59786
rect 455524 59758 455774 59786
rect 455892 59758 456674 59786
rect 456812 59758 457594 59786
rect 458284 59758 458494 59786
rect 458652 59758 459394 59786
rect 459572 59758 460294 59786
rect 460952 59758 461194 59786
rect 461320 59758 462094 59786
rect 462332 59758 462994 59786
rect 463792 59832 463844 59838
rect 463792 59774 463844 59780
rect 463886 59786 463914 60044
rect 464786 59838 464814 60044
rect 464774 59832 464826 59838
rect 452764 22846 452792 59758
rect 452752 22840 452804 22846
rect 452752 22782 452804 22788
rect 454052 20058 454080 59758
rect 455328 57384 455380 57390
rect 455328 57326 455380 57332
rect 454040 20052 454092 20058
rect 454040 19994 454092 20000
rect 452660 14884 452712 14890
rect 452660 14826 452712 14832
rect 453304 9444 453356 9450
rect 453304 9386 453356 9392
rect 450544 8152 450596 8158
rect 450544 8094 450596 8100
rect 452108 8084 452160 8090
rect 452108 8026 452160 8032
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 450924 480 450952 2790
rect 452120 480 452148 8026
rect 453316 480 453344 9386
rect 455340 3738 455368 57326
rect 454500 3732 454552 3738
rect 454500 3674 454552 3680
rect 455328 3732 455380 3738
rect 455328 3674 455380 3680
rect 454512 480 454540 3674
rect 455524 3369 455552 59758
rect 455892 45554 455920 59758
rect 455616 45526 455920 45554
rect 455616 3505 455644 45526
rect 455696 8016 455748 8022
rect 455696 7958 455748 7964
rect 455602 3496 455658 3505
rect 455602 3431 455658 3440
rect 455510 3360 455566 3369
rect 455510 3295 455566 3304
rect 455708 480 455736 7958
rect 456812 3641 456840 59758
rect 458088 57724 458140 57730
rect 458088 57666 458140 57672
rect 456892 9376 456944 9382
rect 456892 9318 456944 9324
rect 456798 3632 456854 3641
rect 456798 3567 456854 3576
rect 456904 480 456932 9318
rect 458100 480 458128 57666
rect 458284 3777 458312 59758
rect 458652 45554 458680 59758
rect 458376 45526 458680 45554
rect 458376 3874 458404 45526
rect 459192 7948 459244 7954
rect 459192 7890 459244 7896
rect 458364 3868 458416 3874
rect 458364 3810 458416 3816
rect 458270 3768 458326 3777
rect 458270 3703 458326 3712
rect 459204 480 459232 7890
rect 459572 3738 459600 59758
rect 460388 9308 460440 9314
rect 460388 9250 460440 9256
rect 459560 3732 459612 3738
rect 459560 3674 459612 3680
rect 460400 480 460428 9250
rect 460952 3942 460980 59758
rect 461320 45554 461348 59758
rect 462228 57180 462280 57186
rect 462228 57122 462280 57128
rect 461044 45526 461348 45554
rect 461044 4010 461072 45526
rect 461032 4004 461084 4010
rect 461032 3946 461084 3952
rect 460940 3936 460992 3942
rect 460940 3878 460992 3884
rect 462240 3534 462268 57122
rect 462332 4078 462360 59758
rect 462780 7880 462832 7886
rect 462780 7822 462832 7828
rect 462320 4072 462372 4078
rect 462320 4014 462372 4020
rect 461584 3528 461636 3534
rect 461584 3470 461636 3476
rect 462228 3528 462280 3534
rect 462228 3470 462280 3476
rect 461596 480 461624 3470
rect 462792 480 462820 7822
rect 463804 3398 463832 59774
rect 463886 59758 463924 59786
rect 465686 59786 465714 60044
rect 464774 59774 464826 59780
rect 463896 4146 463924 59758
rect 465276 59758 465714 59786
rect 466586 59786 466614 60044
rect 467486 59786 467514 60044
rect 466586 59758 466684 59786
rect 463976 9240 464028 9246
rect 463976 9182 464028 9188
rect 463884 4140 463936 4146
rect 463884 4082 463936 4088
rect 463792 3392 463844 3398
rect 463792 3334 463844 3340
rect 463988 480 464016 9182
rect 465172 3528 465224 3534
rect 465172 3470 465224 3476
rect 465184 480 465212 3470
rect 465276 3330 465304 59758
rect 466368 57928 466420 57934
rect 466368 57870 466420 57876
rect 466276 7812 466328 7818
rect 466276 7754 466328 7760
rect 465264 3324 465316 3330
rect 465264 3266 465316 3272
rect 466288 480 466316 7754
rect 466380 3534 466408 57870
rect 466552 57520 466604 57526
rect 466552 57462 466604 57468
rect 466368 3528 466420 3534
rect 466368 3470 466420 3476
rect 466564 3194 466592 57462
rect 466656 3262 466684 59758
rect 467484 59758 467514 59786
rect 468386 59786 468414 60044
rect 469306 59786 469334 60044
rect 470206 59786 470234 60044
rect 471106 59786 471134 60044
rect 468386 59758 468432 59786
rect 469306 59758 469352 59786
rect 467484 57526 467512 59758
rect 468404 57798 468432 59758
rect 468392 57792 468444 57798
rect 468392 57734 468444 57740
rect 467472 57520 467524 57526
rect 467472 57462 467524 57468
rect 469128 57520 469180 57526
rect 469128 57462 469180 57468
rect 468484 16244 468536 16250
rect 468484 16186 468536 16192
rect 467472 9172 467524 9178
rect 467472 9114 467524 9120
rect 466644 3256 466696 3262
rect 466644 3198 466696 3204
rect 466552 3188 466604 3194
rect 466552 3130 466604 3136
rect 467484 480 467512 9114
rect 468496 3806 468524 16186
rect 468484 3800 468536 3806
rect 468484 3742 468536 3748
rect 469140 3534 469168 57462
rect 469324 3670 469352 59758
rect 469416 59758 470234 59786
rect 470612 59758 471134 59786
rect 472006 59786 472034 60044
rect 472906 59786 472934 60044
rect 473806 59786 473834 60044
rect 474706 59786 474734 60044
rect 475626 59786 475654 60044
rect 472006 59758 472112 59786
rect 472906 59758 472940 59786
rect 473806 59758 473860 59786
rect 474706 59758 474872 59786
rect 469312 3664 469364 3670
rect 469312 3606 469364 3612
rect 468668 3528 468720 3534
rect 468668 3470 468720 3476
rect 469128 3528 469180 3534
rect 469128 3470 469180 3476
rect 468680 480 468708 3470
rect 469416 3466 469444 59758
rect 469864 7744 469916 7750
rect 469864 7686 469916 7692
rect 469404 3460 469456 3466
rect 469404 3402 469456 3408
rect 469876 480 469904 7686
rect 470612 3602 470640 59758
rect 471980 57656 472032 57662
rect 471980 57598 472032 57604
rect 471244 13592 471296 13598
rect 471244 13534 471296 13540
rect 471060 9104 471112 9110
rect 471060 9046 471112 9052
rect 470600 3596 470652 3602
rect 470600 3538 470652 3544
rect 471072 480 471100 9046
rect 471256 3466 471284 13534
rect 471992 3738 472020 57598
rect 472084 3874 472112 59758
rect 472912 57662 472940 59758
rect 472900 57656 472952 57662
rect 472900 57598 472952 57604
rect 473832 57458 473860 59758
rect 473820 57452 473872 57458
rect 473820 57394 473872 57400
rect 473268 57180 473320 57186
rect 473268 57122 473320 57128
rect 472072 3868 472124 3874
rect 472072 3810 472124 3816
rect 471980 3732 472032 3738
rect 471980 3674 472032 3680
rect 473280 3534 473308 57122
rect 474556 9036 474608 9042
rect 474556 8978 474608 8984
rect 473452 7676 473504 7682
rect 473452 7618 473504 7624
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 473268 3528 473320 3534
rect 473268 3470 473320 3476
rect 471244 3460 471296 3466
rect 471244 3402 471296 3408
rect 472268 480 472296 3470
rect 473464 480 473492 7618
rect 474568 480 474596 8978
rect 474844 3126 474872 59758
rect 475580 59758 475654 59786
rect 476212 59832 476264 59838
rect 476526 59786 476554 60044
rect 477426 59838 477454 60044
rect 476212 59774 476264 59780
rect 475580 57594 475608 59758
rect 475568 57588 475620 57594
rect 475568 57530 475620 57536
rect 476028 57452 476080 57458
rect 476028 57394 476080 57400
rect 476040 6914 476068 57394
rect 475764 6886 476068 6914
rect 474832 3120 474884 3126
rect 474832 3062 474884 3068
rect 475764 480 475792 6886
rect 476224 2990 476252 59774
rect 476316 59758 476554 59786
rect 477414 59832 477466 59838
rect 477414 59774 477466 59780
rect 478326 59786 478354 60044
rect 479226 59786 479254 60044
rect 480126 59786 480154 60044
rect 481026 59786 481054 60044
rect 481946 59786 481974 60044
rect 478326 59758 478368 59786
rect 476316 3058 476344 59758
rect 478340 57866 478368 59758
rect 478984 59758 479254 59786
rect 480088 59758 480154 59786
rect 480272 59758 481054 59786
rect 481928 59758 481974 59786
rect 482846 59786 482874 60044
rect 483746 59786 483774 60044
rect 484646 59786 484674 60044
rect 485546 59786 485574 60044
rect 486446 59786 486474 60044
rect 487366 59786 487394 60044
rect 482846 59758 482876 59786
rect 483746 59758 483796 59786
rect 478328 57860 478380 57866
rect 478328 57802 478380 57808
rect 478144 8968 478196 8974
rect 478144 8910 478196 8916
rect 476948 7608 477000 7614
rect 476948 7550 477000 7556
rect 476304 3052 476356 3058
rect 476304 2994 476356 3000
rect 476212 2984 476264 2990
rect 476212 2926 476264 2932
rect 476960 480 476988 7550
rect 478156 480 478184 8910
rect 478984 2922 479012 59758
rect 480088 57118 480116 59758
rect 480168 57656 480220 57662
rect 480168 57598 480220 57604
rect 480076 57112 480128 57118
rect 480076 57054 480128 57060
rect 480180 3534 480208 57598
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 478972 2916 479024 2922
rect 478972 2858 479024 2864
rect 479352 480 479380 3470
rect 480272 2854 480300 59758
rect 481928 57390 481956 59758
rect 482848 57730 482876 59758
rect 483768 57798 483796 59758
rect 484596 59758 484674 59786
rect 485516 59758 485574 59786
rect 486436 59758 486474 59786
rect 487356 59758 487394 59786
rect 488266 59786 488294 60044
rect 489166 59786 489194 60044
rect 490066 59922 490094 60044
rect 490024 59894 490094 59922
rect 488266 59758 488304 59786
rect 489166 59758 489224 59786
rect 484596 57934 484624 59758
rect 484584 57928 484636 57934
rect 484584 57870 484636 57876
rect 483756 57792 483808 57798
rect 483756 57734 483808 57740
rect 482836 57724 482888 57730
rect 482836 57666 482888 57672
rect 482928 57588 482980 57594
rect 482928 57530 482980 57536
rect 481916 57384 481968 57390
rect 481916 57326 481968 57332
rect 481640 29640 481692 29646
rect 481640 29582 481692 29588
rect 481652 16574 481680 29582
rect 481652 16546 481772 16574
rect 480536 8152 480588 8158
rect 480536 8094 480588 8100
rect 480260 2848 480312 2854
rect 480260 2790 480312 2796
rect 480548 480 480576 8094
rect 481744 480 481772 16546
rect 482940 6914 482968 57530
rect 485516 57526 485544 59758
rect 485504 57520 485556 57526
rect 485504 57462 485556 57468
rect 486436 57186 486464 59758
rect 487356 57458 487384 59758
rect 488276 57662 488304 59758
rect 488264 57656 488316 57662
rect 488264 57598 488316 57604
rect 489196 57594 489224 59758
rect 489184 57588 489236 57594
rect 489184 57530 489236 57536
rect 487344 57452 487396 57458
rect 487344 57394 487396 57400
rect 489184 57316 489236 57322
rect 489184 57258 489236 57264
rect 486424 57180 486476 57186
rect 486424 57122 486476 57128
rect 487068 56636 487120 56642
rect 487068 56578 487120 56584
rect 483664 55956 483716 55962
rect 483664 55898 483716 55904
rect 483676 16574 483704 55898
rect 485044 55888 485096 55894
rect 485044 55830 485096 55836
rect 483676 16546 483796 16574
rect 483664 14476 483716 14482
rect 483664 14418 483716 14424
rect 482848 6886 482968 6914
rect 482848 480 482876 6886
rect 483676 3482 483704 14418
rect 483768 3602 483796 16546
rect 484768 12232 484820 12238
rect 484768 12174 484820 12180
rect 483756 3596 483808 3602
rect 483756 3538 483808 3544
rect 483676 3454 484072 3482
rect 484044 480 484072 3454
rect 484780 490 484808 12174
rect 485056 3126 485084 55830
rect 486424 25560 486476 25566
rect 486424 25502 486476 25508
rect 486436 3670 486464 25502
rect 486424 3664 486476 3670
rect 486424 3606 486476 3612
rect 487080 3534 487108 56578
rect 489196 3670 489224 57258
rect 490024 56642 490052 59894
rect 490966 59786 490994 60044
rect 491866 59786 491894 60044
rect 490116 59758 490994 59786
rect 491864 59758 491894 59786
rect 492766 59786 492794 60044
rect 493686 59786 493714 60044
rect 494586 59786 494614 60044
rect 495486 59786 495514 60044
rect 496386 59786 496414 60044
rect 497286 59786 497314 60044
rect 498186 59786 498214 60044
rect 499086 59786 499114 60044
rect 500006 59786 500034 60044
rect 500906 59786 500934 60044
rect 501806 59786 501834 60044
rect 492766 59758 492812 59786
rect 493686 59758 494008 59786
rect 494586 59758 494652 59786
rect 495486 59758 495572 59786
rect 496386 59758 496676 59786
rect 497286 59758 497320 59786
rect 498186 59758 498240 59786
rect 499086 59758 499528 59786
rect 500006 59758 500080 59786
rect 490012 56636 490064 56642
rect 490012 56578 490064 56584
rect 489276 11892 489328 11898
rect 489276 11834 489328 11840
rect 489288 4146 489316 11834
rect 490116 6914 490144 59758
rect 491864 57662 491892 59758
rect 491852 57656 491904 57662
rect 491852 57598 491904 57604
rect 492784 57594 492812 59758
rect 492864 57656 492916 57662
rect 492864 57598 492916 57604
rect 492772 57588 492824 57594
rect 492772 57530 492824 57536
rect 492876 16574 492904 57598
rect 493876 57588 493928 57594
rect 493876 57530 493928 57536
rect 492876 16546 493088 16574
rect 490564 12096 490616 12102
rect 490564 12038 490616 12044
rect 489932 6886 490144 6914
rect 489276 4140 489328 4146
rect 489276 4082 489328 4088
rect 488816 3664 488868 3670
rect 488816 3606 488868 3612
rect 489184 3664 489236 3670
rect 489184 3606 489236 3612
rect 486424 3528 486476 3534
rect 486424 3470 486476 3476
rect 487068 3528 487120 3534
rect 487068 3470 487120 3476
rect 485044 3120 485096 3126
rect 485044 3062 485096 3068
rect 485056 598 485268 626
rect 485056 490 485084 598
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 462 485084 490
rect 485240 480 485268 598
rect 486436 480 486464 3470
rect 487620 3120 487672 3126
rect 487620 3062 487672 3068
rect 487632 480 487660 3062
rect 488828 480 488856 3606
rect 489932 480 489960 6886
rect 490576 2990 490604 12038
rect 491116 4140 491168 4146
rect 491116 4082 491168 4088
rect 490564 2984 490616 2990
rect 490564 2926 490616 2932
rect 491128 480 491156 4082
rect 492312 2984 492364 2990
rect 492312 2926 492364 2932
rect 492324 480 492352 2926
rect 493060 490 493088 16546
rect 493888 3194 493916 57530
rect 493980 3398 494008 59758
rect 494624 57662 494652 59758
rect 495544 57662 495572 59758
rect 494612 57656 494664 57662
rect 494612 57598 494664 57604
rect 495348 57656 495400 57662
rect 495348 57598 495400 57604
rect 495532 57656 495584 57662
rect 495532 57598 495584 57604
rect 495360 3874 495388 57598
rect 495348 3868 495400 3874
rect 495348 3810 495400 3816
rect 496648 3806 496676 59758
rect 497292 57662 497320 59758
rect 498212 57662 498240 59758
rect 496728 57656 496780 57662
rect 496728 57598 496780 57604
rect 497280 57656 497332 57662
rect 497280 57598 497332 57604
rect 498108 57656 498160 57662
rect 498108 57598 498160 57604
rect 498200 57656 498252 57662
rect 498200 57598 498252 57604
rect 499396 57656 499448 57662
rect 499396 57598 499448 57604
rect 495900 3800 495952 3806
rect 495900 3742 495952 3748
rect 496636 3800 496688 3806
rect 496636 3742 496688 3748
rect 494704 3664 494756 3670
rect 494704 3606 494756 3612
rect 493968 3392 494020 3398
rect 493968 3334 494020 3340
rect 493876 3188 493928 3194
rect 493876 3130 493928 3136
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 3606
rect 495912 480 495940 3742
rect 496740 3738 496768 57598
rect 497464 13388 497516 13394
rect 497464 13330 497516 13336
rect 496728 3732 496780 3738
rect 496728 3674 496780 3680
rect 497096 3188 497148 3194
rect 497096 3130 497148 3136
rect 497108 480 497136 3130
rect 497476 3058 497504 13330
rect 498120 3670 498148 57598
rect 499408 6914 499436 57598
rect 499316 6886 499436 6914
rect 498108 3664 498160 3670
rect 498108 3606 498160 3612
rect 498200 3596 498252 3602
rect 498200 3538 498252 3544
rect 497464 3052 497516 3058
rect 497464 2994 497516 3000
rect 498212 480 498240 3538
rect 499316 2854 499344 6886
rect 499396 3052 499448 3058
rect 499396 2994 499448 3000
rect 499304 2848 499356 2854
rect 499304 2790 499356 2796
rect 499408 480 499436 2994
rect 499500 2922 499528 59758
rect 500052 57662 500080 59758
rect 500880 59758 500934 59786
rect 501800 59758 501834 59786
rect 502706 59786 502734 60044
rect 503606 59786 503634 60044
rect 504506 59786 504534 60044
rect 505426 59786 505454 60044
rect 506326 59786 506354 60044
rect 502706 59758 502748 59786
rect 503606 59758 503668 59786
rect 504506 59758 504588 59786
rect 505426 59758 505508 59786
rect 500040 57656 500092 57662
rect 500040 57598 500092 57604
rect 500776 57656 500828 57662
rect 500776 57598 500828 57604
rect 500592 3392 500644 3398
rect 500592 3334 500644 3340
rect 499488 2916 499540 2922
rect 499488 2858 499540 2864
rect 500604 480 500632 3334
rect 500788 2990 500816 57598
rect 500880 3058 500908 59758
rect 501800 57662 501828 59758
rect 501788 57656 501840 57662
rect 501788 57598 501840 57604
rect 502248 57656 502300 57662
rect 502248 57598 502300 57604
rect 501604 56228 501656 56234
rect 501604 56170 501656 56176
rect 501328 11824 501380 11830
rect 501328 11766 501380 11772
rect 500868 3052 500920 3058
rect 500868 2994 500920 3000
rect 500776 2984 500828 2990
rect 500776 2926 500828 2932
rect 501340 490 501368 11766
rect 501616 3534 501644 56170
rect 501604 3528 501656 3534
rect 501604 3470 501656 3476
rect 502260 3126 502288 57598
rect 502720 57050 502748 59758
rect 502708 57044 502760 57050
rect 502708 56986 502760 56992
rect 503536 57044 503588 57050
rect 503536 56986 503588 56992
rect 502984 3460 503036 3466
rect 502984 3402 503036 3408
rect 502248 3120 502300 3126
rect 502248 3062 502300 3068
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 3402
rect 503548 3194 503576 56986
rect 503640 3262 503668 59758
rect 504560 57186 504588 59758
rect 505480 57662 505508 59758
rect 506308 59758 506354 59786
rect 507226 59786 507254 60044
rect 508126 59786 508154 60044
rect 509026 59786 509054 60044
rect 509926 59786 509954 60044
rect 510826 59786 510854 60044
rect 507226 59758 507256 59786
rect 508126 59758 508176 59786
rect 509026 59758 509188 59786
rect 505468 57656 505520 57662
rect 505468 57598 505520 57604
rect 504548 57180 504600 57186
rect 504548 57122 504600 57128
rect 505008 57180 505060 57186
rect 505008 57122 505060 57128
rect 504364 13116 504416 13122
rect 504364 13058 504416 13064
rect 504180 3868 504232 3874
rect 504180 3810 504232 3816
rect 503628 3256 503680 3262
rect 503628 3198 503680 3204
rect 503536 3188 503588 3194
rect 503536 3130 503588 3136
rect 504192 480 504220 3810
rect 504376 3534 504404 13058
rect 504364 3528 504416 3534
rect 504364 3470 504416 3476
rect 505020 3330 505048 57122
rect 506308 4146 506336 59758
rect 507228 57662 507256 59758
rect 508148 57662 508176 59758
rect 506388 57656 506440 57662
rect 506388 57598 506440 57604
rect 507216 57656 507268 57662
rect 507216 57598 507268 57604
rect 507768 57656 507820 57662
rect 507768 57598 507820 57604
rect 508136 57656 508188 57662
rect 508136 57598 508188 57604
rect 509056 57656 509108 57662
rect 509056 57598 509108 57604
rect 506296 4140 506348 4146
rect 506296 4082 506348 4088
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 505008 3324 505060 3330
rect 505008 3266 505060 3272
rect 505388 480 505416 3470
rect 506400 3398 506428 57598
rect 507124 57248 507176 57254
rect 507124 57190 507176 57196
rect 506480 10328 506532 10334
rect 506480 10270 506532 10276
rect 506388 3392 506440 3398
rect 506388 3334 506440 3340
rect 506492 480 506520 10270
rect 507136 3534 507164 57190
rect 507780 4078 507808 57598
rect 507768 4072 507820 4078
rect 507768 4014 507820 4020
rect 509068 4010 509096 57598
rect 509056 4004 509108 4010
rect 509056 3946 509108 3952
rect 509160 3942 509188 59758
rect 509896 59758 509954 59786
rect 510816 59758 510854 59786
rect 511746 59786 511774 60044
rect 512646 59786 512674 60044
rect 513546 59786 513574 60044
rect 514446 59786 514474 60044
rect 515346 59786 515374 60044
rect 516246 59786 516274 60044
rect 511746 59758 511948 59786
rect 512646 59758 512684 59786
rect 513546 59758 513604 59786
rect 514446 59758 514708 59786
rect 509896 57662 509924 59758
rect 510816 57662 510844 59758
rect 509884 57656 509936 57662
rect 509884 57598 509936 57604
rect 510528 57656 510580 57662
rect 510528 57598 510580 57604
rect 510804 57656 510856 57662
rect 510804 57598 510856 57604
rect 511816 57656 511868 57662
rect 511816 57598 511868 57604
rect 509148 3936 509200 3942
rect 509148 3878 509200 3884
rect 510540 3874 510568 57598
rect 510528 3868 510580 3874
rect 510528 3810 510580 3816
rect 511828 3806 511856 57598
rect 511816 3800 511868 3806
rect 511816 3742 511868 3748
rect 511920 3738 511948 59758
rect 512656 57458 512684 59758
rect 513576 57662 513604 59758
rect 513564 57656 513616 57662
rect 513564 57598 513616 57604
rect 514576 57656 514628 57662
rect 514576 57598 514628 57604
rect 512644 57452 512696 57458
rect 512644 57394 512696 57400
rect 513288 57452 513340 57458
rect 513288 57394 513340 57400
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 507676 3732 507728 3738
rect 507676 3674 507728 3680
rect 511908 3732 511960 3738
rect 511908 3674 511960 3680
rect 507124 3528 507176 3534
rect 507124 3470 507176 3476
rect 507688 480 507716 3674
rect 511264 3664 511316 3670
rect 511264 3606 511316 3612
rect 508872 3528 508924 3534
rect 508872 3470 508924 3476
rect 508884 480 508912 3470
rect 510068 3460 510120 3466
rect 510068 3402 510120 3408
rect 510080 480 510108 3402
rect 511276 480 511304 3606
rect 512472 480 512500 4218
rect 513300 3670 513328 57394
rect 513564 5636 513616 5642
rect 513564 5578 513616 5584
rect 513288 3664 513340 3670
rect 513288 3606 513340 3612
rect 513576 480 513604 5578
rect 514588 3534 514616 57598
rect 514576 3528 514628 3534
rect 514576 3470 514628 3476
rect 514680 3466 514708 59758
rect 515324 59758 515374 59786
rect 516244 59758 516274 59786
rect 516846 59786 516874 60044
rect 516846 59758 516916 59786
rect 515324 57662 515352 59758
rect 515312 57656 515364 57662
rect 515312 57598 515364 57604
rect 516048 57656 516100 57662
rect 516048 57598 516100 57604
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 514760 3596 514812 3602
rect 514760 3538 514812 3544
rect 514668 3460 514720 3466
rect 514668 3402 514720 3408
rect 514772 480 514800 3538
rect 515968 480 515996 4286
rect 516060 3505 516088 57598
rect 516244 57594 516272 59758
rect 516888 57662 516916 59758
rect 516876 57656 516928 57662
rect 516876 57598 516928 57604
rect 517428 57656 517480 57662
rect 517428 57598 517480 57604
rect 516232 57588 516284 57594
rect 516232 57530 516284 57536
rect 517336 57588 517388 57594
rect 517336 57530 517388 57536
rect 517152 5704 517204 5710
rect 517152 5646 517204 5652
rect 516046 3496 516102 3505
rect 516046 3431 516102 3440
rect 517164 480 517192 5646
rect 517348 3602 517376 57530
rect 517336 3596 517388 3602
rect 517336 3538 517388 3544
rect 517440 3369 517468 57598
rect 519556 6866 519584 60415
rect 519648 20670 519676 71023
rect 519740 33114 519768 82175
rect 519832 46918 519860 93191
rect 519924 60722 519952 104343
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 519912 60716 519964 60722
rect 519912 60658 519964 60664
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 519820 46912 519872 46918
rect 519820 46854 519872 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 519728 33108 519780 33114
rect 580170 33079 580172 33088
rect 519728 33050 519780 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 519636 20664 519688 20670
rect 519636 20606 519688 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 519544 6860 519596 6866
rect 519544 6802 519596 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 545488 6792 545540 6798
rect 545488 6734 545540 6740
rect 538404 6112 538456 6118
rect 538404 6054 538456 6060
rect 534908 6044 534960 6050
rect 534908 5986 534960 5992
rect 531320 5976 531372 5982
rect 531320 5918 531372 5924
rect 527824 5908 527876 5914
rect 527824 5850 527876 5856
rect 524236 5840 524288 5846
rect 524236 5782 524288 5788
rect 520740 5772 520792 5778
rect 520740 5714 520792 5720
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 517426 3360 517482 3369
rect 517426 3295 517482 3304
rect 518348 2848 518400 2854
rect 518348 2790 518400 2796
rect 518360 480 518388 2790
rect 519556 480 519584 4354
rect 520752 480 520780 5714
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 521844 2916 521896 2922
rect 521844 2858 521896 2864
rect 521856 480 521884 2858
rect 523052 480 523080 4422
rect 524248 480 524276 5782
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 525432 2984 525484 2990
rect 525432 2926 525484 2932
rect 525444 480 525472 2926
rect 526640 480 526668 4490
rect 527836 480 527864 5850
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 529020 3052 529072 3058
rect 529020 2994 529072 3000
rect 529032 480 529060 2994
rect 530136 480 530164 4558
rect 531332 480 531360 5918
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 3120 532568 3126
rect 532516 3062 532568 3068
rect 532528 480 532556 3062
rect 533724 480 533752 4626
rect 534920 480 534948 5986
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 536104 3188 536156 3194
rect 536104 3130 536156 3136
rect 536116 480 536144 3130
rect 537220 480 537248 4694
rect 538416 480 538444 6054
rect 541992 5568 542044 5574
rect 541992 5510 542044 5516
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3256 539652 3262
rect 539600 3198 539652 3204
rect 539612 480 539640 3198
rect 540808 480 540836 5442
rect 542004 480 542032 5510
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 3324 543240 3330
rect 543188 3266 543240 3272
rect 543200 480 543228 3266
rect 544396 480 544424 5374
rect 545500 480 545528 6734
rect 549076 6724 549128 6730
rect 549076 6666 549128 6672
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 3392 546736 3398
rect 546684 3334 546736 3340
rect 546696 480 546724 3334
rect 547892 480 547920 5306
rect 549088 480 549116 6666
rect 552664 6656 552716 6662
rect 580184 6633 580212 6802
rect 552664 6598 552716 6604
rect 580170 6624 580226 6633
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 4140 550324 4146
rect 550272 4082 550324 4088
rect 550284 480 550312 4082
rect 551480 480 551508 5238
rect 552676 480 552704 6598
rect 556160 6588 556212 6594
rect 580170 6559 580226 6568
rect 556160 6530 556212 6536
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 4072 553820 4078
rect 553768 4014 553820 4020
rect 553780 480 553808 4014
rect 554976 480 555004 5170
rect 556172 480 556200 6530
rect 559748 6520 559800 6526
rect 559748 6462 559800 6468
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 4004 557408 4010
rect 557356 3946 557408 3952
rect 557368 480 557396 3946
rect 558564 480 558592 5102
rect 559760 480 559788 6462
rect 563244 6452 563296 6458
rect 563244 6394 563296 6400
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560852 3936 560904 3942
rect 560852 3878 560904 3884
rect 560864 480 560892 3878
rect 562060 480 562088 5034
rect 563256 480 563284 6394
rect 566832 6384 566884 6390
rect 566832 6326 566884 6332
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3868 564492 3874
rect 564440 3810 564492 3816
rect 564452 480 564480 3810
rect 565648 480 565676 4966
rect 566844 480 566872 6326
rect 570328 6316 570380 6322
rect 570328 6258 570380 6264
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3800 568080 3806
rect 568028 3742 568080 3748
rect 568040 480 568068 3742
rect 569144 480 569172 4898
rect 570340 480 570368 6258
rect 573916 6248 573968 6254
rect 573916 6190 573968 6196
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3732 571576 3738
rect 571524 3674 571576 3680
rect 571536 480 571564 3674
rect 572732 480 572760 4830
rect 573928 480 573956 6190
rect 577412 6180 577464 6186
rect 577412 6122 577464 6128
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3664 575164 3670
rect 575112 3606 575164 3612
rect 575124 480 575152 3606
rect 576320 480 576348 4762
rect 577424 480 577452 6122
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 580998 3496 581054 3505
rect 578620 480 578648 3470
rect 579804 3460 579856 3466
rect 580998 3431 581054 3440
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3431
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 684256 3570 684312
rect 3422 632032 3478 632088
rect 3606 671200 3662 671256
rect 3514 619112 3570 619168
rect 3422 579944 3478 580000
rect 3698 658144 3754 658200
rect 3606 606056 3662 606112
rect 3514 566888 3570 566944
rect 3790 645088 3846 645144
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 519542 636792 519598 636848
rect 69018 636656 69074 636712
rect 69018 626320 69074 626376
rect 69018 615460 69074 615496
rect 69018 615440 69020 615460
rect 69020 615440 69072 615460
rect 69072 615440 69074 615460
rect 69018 604560 69074 604616
rect 69018 593680 69074 593736
rect 3698 593000 3754 593056
rect 3606 553832 3662 553888
rect 3422 527856 3478 527912
rect 69018 582800 69074 582856
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 519634 626184 519690 626240
rect 519542 581712 519598 581768
rect 69018 571920 69074 571976
rect 69018 560904 69074 560960
rect 69018 550160 69074 550216
rect 3698 540776 3754 540832
rect 3514 514800 3570 514856
rect 3422 488688 3478 488744
rect 69018 539144 69074 539200
rect 580170 670656 580226 670692
rect 580170 657328 580226 657384
rect 519726 615032 519782 615088
rect 580170 644000 580226 644056
rect 519818 603880 519874 603936
rect 519634 570560 519690 570616
rect 519542 537376 519598 537432
rect 69018 528264 69074 528320
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580170 604152 580226 604208
rect 519910 592864 519966 592920
rect 579802 590960 579858 591016
rect 519726 559544 519782 559600
rect 519634 526224 519690 526280
rect 69018 517420 69020 517440
rect 69020 517420 69072 517440
rect 69072 517420 69074 517440
rect 69018 517384 69074 517420
rect 69018 506504 69074 506560
rect 3606 501744 3662 501800
rect 3514 475632 3570 475688
rect 69018 495624 69074 495680
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 551112 580226 551168
rect 519818 548392 519874 548448
rect 580170 537784 580226 537840
rect 519726 515072 519782 515128
rect 519542 492768 519598 492824
rect 69018 484744 69074 484800
rect 69018 473864 69074 473920
rect 69018 462984 69074 463040
rect 3606 462576 3662 462632
rect 3422 449520 3478 449576
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 519818 504056 519874 504112
rect 580170 497936 580226 497992
rect 519634 481752 519690 481808
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 519726 470736 519782 470792
rect 519542 459584 519598 459640
rect 69018 452104 69074 452160
rect 69018 441224 69074 441280
rect 580170 458088 580226 458144
rect 519634 448568 519690 448624
rect 580170 444760 580226 444816
rect 519542 437416 519598 437472
rect 3514 436600 3570 436656
rect 3422 423544 3478 423600
rect 69018 430344 69074 430400
rect 69018 419328 69074 419384
rect 580170 431568 580226 431624
rect 519634 426264 519690 426320
rect 580170 418240 580226 418296
rect 519542 415248 519598 415304
rect 3514 410488 3570 410544
rect 69018 408584 69074 408640
rect 69018 397568 69074 397624
rect 3422 397432 3478 397488
rect 580170 404912 580226 404968
rect 519634 404096 519690 404152
rect 519542 392944 519598 393000
rect 580170 391720 580226 391776
rect 69018 386688 69074 386744
rect 3422 384376 3478 384432
rect 519542 381928 519598 381984
rect 580170 378392 580226 378448
rect 69018 375808 69074 375864
rect 3422 371320 3478 371376
rect 519542 370776 519598 370832
rect 580170 365064 580226 365120
rect 69018 364928 69074 364984
rect 519358 359760 519414 359816
rect 3422 358400 3478 358456
rect 69018 354048 69074 354104
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 519818 348608 519874 348664
rect 3146 345344 3202 345400
rect 69018 343168 69074 343224
rect 580170 338544 580226 338600
rect 520002 337456 520058 337512
rect 3422 332288 3478 332344
rect 69018 332152 69074 332208
rect 519358 326304 519414 326360
rect 580170 325216 580226 325272
rect 69018 321272 69074 321328
rect 3422 319232 3478 319288
rect 520186 315288 520242 315344
rect 580170 312024 580226 312080
rect 69018 310392 69074 310448
rect 3422 306176 3478 306232
rect 519358 304136 519414 304192
rect 69018 299532 69074 299568
rect 69018 299512 69020 299532
rect 69020 299512 69072 299532
rect 69072 299512 69074 299532
rect 580170 298696 580226 298752
rect 3422 293120 3478 293176
rect 519542 293120 519598 293176
rect 69018 288632 69074 288688
rect 580170 285368 580226 285424
rect 519542 281968 519598 282024
rect 3422 280064 3478 280120
rect 69018 277752 69074 277808
rect 580170 272176 580226 272232
rect 519542 270816 519598 270872
rect 3514 267144 3570 267200
rect 69018 266872 69074 266928
rect 519634 259800 519690 259856
rect 69018 255992 69074 256048
rect 3422 254088 3478 254144
rect 519542 248648 519598 248704
rect 69018 245112 69074 245168
rect 3514 241032 3570 241088
rect 69018 234232 69074 234288
rect 3422 227976 3478 228032
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 519634 237496 519690 237552
rect 519542 226480 519598 226536
rect 69018 223352 69074 223408
rect 3514 214920 3570 214976
rect 69018 212472 69074 212528
rect 3422 201864 3478 201920
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 519726 215328 519782 215384
rect 519634 204312 519690 204368
rect 69018 201592 69074 201648
rect 519542 193160 519598 193216
rect 69018 190576 69074 190632
rect 3606 188808 3662 188864
rect 69018 179696 69074 179752
rect 3514 175888 3570 175944
rect 3422 162832 3478 162888
rect 69018 168816 69074 168872
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 519726 182008 519782 182064
rect 519634 170992 519690 171048
rect 519542 159840 519598 159896
rect 69018 157936 69074 157992
rect 3606 149776 3662 149832
rect 69018 147056 69074 147112
rect 3514 136720 3570 136776
rect 3422 123664 3478 123720
rect 69018 136176 69074 136232
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 519818 148688 519874 148744
rect 519726 137672 519782 137728
rect 519634 126520 519690 126576
rect 69018 125296 69074 125352
rect 519542 115504 519598 115560
rect 69018 114416 69074 114472
rect 3698 110608 3754 110664
rect 69018 103556 69074 103592
rect 69018 103536 69020 103556
rect 69020 103536 69072 103556
rect 69072 103536 69074 103556
rect 3606 97552 3662 97608
rect 3514 84632 3570 84688
rect 3422 71576 3478 71632
rect 69018 92656 69074 92712
rect 69018 81776 69074 81832
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 519910 104352 519966 104408
rect 519818 93200 519874 93256
rect 519726 82184 519782 82240
rect 519634 71032 519690 71088
rect 69018 70760 69074 70816
rect 519542 60424 519598 60480
rect 69018 60152 69074 60208
rect 3790 58520 3846 58576
rect 3698 45464 3754 45520
rect 3606 32408 3662 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 11150 3440 11206 3496
rect 19430 3712 19486 3768
rect 20626 3576 20682 3632
rect 133970 3712 134026 3768
rect 161570 3440 161626 3496
rect 162950 3576 163006 3632
rect 165710 3304 165766 3360
rect 351642 3304 351698 3360
rect 355230 3440 355286 3496
rect 358726 3576 358782 3632
rect 362314 3712 362370 3768
rect 455602 3440 455658 3496
rect 455510 3304 455566 3360
rect 456798 3576 456854 3632
rect 458270 3712 458326 3768
rect 516046 3440 516102 3496
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 517426 3304 517482 3360
rect 580170 6568 580226 6624
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3601 671258 3667 671261
rect -960 671256 3667 671258
rect -960 671200 3606 671256
rect 3662 671200 3667 671256
rect -960 671198 3667 671200
rect -960 671108 480 671198
rect 3601 671195 3667 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3693 658202 3759 658205
rect -960 658200 3759 658202
rect -960 658144 3698 658200
rect 3754 658144 3759 658200
rect -960 658142 3759 658144
rect -960 658052 480 658142
rect 3693 658139 3759 658142
rect 580165 657386 580231 657389
rect 583520 657386 584960 657476
rect 580165 657384 584960 657386
rect 580165 657328 580170 657384
rect 580226 657328 584960 657384
rect 580165 657326 584960 657328
rect 580165 657323 580231 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 3785 645146 3851 645149
rect -960 645144 3851 645146
rect -960 645088 3790 645144
rect 3846 645088 3851 645144
rect -960 645086 3851 645088
rect -960 644996 480 645086
rect 3785 645083 3851 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 519537 636850 519603 636853
rect 517654 636848 519603 636850
rect 517654 636799 519542 636848
rect 517132 636792 519542 636799
rect 519598 636792 519603 636848
rect 517132 636790 519603 636792
rect 517132 636739 517714 636790
rect 519537 636787 519603 636790
rect 69013 636714 69079 636717
rect 69013 636712 71514 636714
rect 69013 636656 69018 636712
rect 69074 636682 71514 636712
rect 69074 636656 72036 636682
rect 69013 636654 72036 636656
rect 69013 636651 69079 636654
rect 71454 636622 72036 636654
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 69013 626378 69079 626381
rect 69013 626376 71514 626378
rect 69013 626320 69018 626376
rect 69074 626352 71514 626376
rect 69074 626320 72036 626352
rect 69013 626318 72036 626320
rect 69013 626315 69079 626318
rect 71454 626292 72036 626318
rect 519629 626242 519695 626245
rect 517654 626240 519695 626242
rect 517654 626184 519634 626240
rect 519690 626184 519695 626240
rect 517654 626182 519695 626184
rect 517654 626156 517714 626182
rect 519629 626179 519695 626182
rect 517132 626096 517714 626156
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 69013 615498 69079 615501
rect 69013 615496 71514 615498
rect 69013 615440 69018 615496
rect 69074 615474 71514 615496
rect 69074 615440 72036 615474
rect 69013 615438 72036 615440
rect 69013 615435 69079 615438
rect 71454 615414 72036 615438
rect 519721 615090 519787 615093
rect 517654 615088 519787 615090
rect 517654 615063 519726 615088
rect 517132 615032 519726 615063
rect 519782 615032 519787 615088
rect 517132 615030 519787 615032
rect 517132 615003 517714 615030
rect 519721 615027 519787 615030
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 69013 604618 69079 604621
rect 69013 604616 71514 604618
rect 69013 604560 69018 604616
rect 69074 604577 71514 604616
rect 69074 604560 72036 604577
rect 69013 604558 72036 604560
rect 69013 604555 69079 604558
rect 71454 604517 72036 604558
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 517132 603938 517714 603950
rect 519813 603938 519879 603941
rect 517132 603936 519879 603938
rect 517132 603890 519818 603936
rect 517654 603880 519818 603890
rect 519874 603880 519879 603936
rect 517654 603878 519879 603880
rect 519813 603875 519879 603878
rect 69013 593738 69079 593741
rect 69013 593736 71514 593738
rect 69013 593680 69018 593736
rect 69074 593680 71514 593736
rect 69013 593679 71514 593680
rect 69013 593678 72036 593679
rect 69013 593675 69079 593678
rect 71454 593619 72036 593678
rect -960 593058 480 593148
rect 3693 593058 3759 593061
rect -960 593056 3759 593058
rect -960 593000 3698 593056
rect 3754 593000 3759 593056
rect -960 592998 3759 593000
rect -960 592908 480 592998
rect 3693 592995 3759 592998
rect 519905 592922 519971 592925
rect 517654 592920 519971 592922
rect 517654 592864 519910 592920
rect 519966 592864 519971 592920
rect 517654 592862 519971 592864
rect 517654 592856 517714 592862
rect 519905 592859 519971 592862
rect 517132 592796 517714 592856
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 69013 582858 69079 582861
rect 69013 582856 71514 582858
rect 69013 582800 69018 582856
rect 69074 582801 71514 582856
rect 69074 582800 72036 582801
rect 69013 582798 72036 582800
rect 69013 582795 69079 582798
rect 71454 582741 72036 582798
rect 519537 581770 519603 581773
rect 517654 581768 519603 581770
rect 517654 581743 519542 581768
rect 517132 581712 519542 581743
rect 519598 581712 519603 581768
rect 517132 581710 519603 581712
rect 517132 581683 517714 581710
rect 519537 581707 519603 581710
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 69013 571978 69079 571981
rect 69013 571976 71514 571978
rect 69013 571920 69018 571976
rect 69074 571920 71514 571976
rect 69013 571918 71514 571920
rect 69013 571915 69079 571918
rect 71454 571904 71514 571918
rect 71454 571844 72036 571904
rect 517132 570618 517714 570649
rect 519629 570618 519695 570621
rect 517132 570616 519695 570618
rect 517132 570589 519634 570616
rect 517654 570560 519634 570589
rect 519690 570560 519695 570616
rect 517654 570558 519695 570560
rect 519629 570555 519695 570558
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 69013 560962 69079 560965
rect 71454 560962 72036 561006
rect 69013 560960 72036 560962
rect 69013 560904 69018 560960
rect 69074 560946 72036 560960
rect 69074 560904 71514 560946
rect 69013 560902 71514 560904
rect 69013 560899 69079 560902
rect 519721 559602 519787 559605
rect 517654 559600 519787 559602
rect 517654 559556 519726 559600
rect 517132 559544 519726 559556
rect 519782 559544 519787 559600
rect 517132 559542 519787 559544
rect 517132 559496 517714 559542
rect 519721 559539 519787 559542
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 580165 551170 580231 551173
rect 583520 551170 584960 551260
rect 580165 551168 584960 551170
rect 580165 551112 580170 551168
rect 580226 551112 584960 551168
rect 580165 551110 584960 551112
rect 580165 551107 580231 551110
rect 583520 551020 584960 551110
rect 69013 550218 69079 550221
rect 69013 550216 71514 550218
rect 69013 550160 69018 550216
rect 69074 550160 71514 550216
rect 69013 550158 71514 550160
rect 69013 550155 69079 550158
rect 71454 550128 71514 550158
rect 71454 550068 72036 550128
rect 519813 548450 519879 548453
rect 517654 548448 519879 548450
rect 517654 548442 519818 548448
rect 517132 548392 519818 548442
rect 519874 548392 519879 548448
rect 517132 548390 519879 548392
rect 517132 548382 517714 548390
rect 519813 548387 519879 548390
rect -960 540834 480 540924
rect 3693 540834 3759 540837
rect -960 540832 3759 540834
rect -960 540776 3698 540832
rect 3754 540776 3759 540832
rect -960 540774 3759 540776
rect -960 540684 480 540774
rect 3693 540771 3759 540774
rect 69013 539202 69079 539205
rect 71454 539202 72036 539230
rect 69013 539200 72036 539202
rect 69013 539144 69018 539200
rect 69074 539170 72036 539200
rect 69074 539144 71514 539170
rect 69013 539142 71514 539144
rect 69013 539139 69079 539142
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 519537 537434 519603 537437
rect 517654 537432 519603 537434
rect 517654 537376 519542 537432
rect 519598 537376 519603 537432
rect 517654 537374 519603 537376
rect 517654 537349 517714 537374
rect 519537 537371 519603 537374
rect 517132 537289 517714 537349
rect 69013 528322 69079 528325
rect 71454 528322 72036 528333
rect 69013 528320 72036 528322
rect 69013 528264 69018 528320
rect 69074 528273 72036 528320
rect 69074 528264 71514 528273
rect 69013 528262 71514 528264
rect 69013 528259 69079 528262
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 519629 526282 519695 526285
rect 517654 526280 519695 526282
rect 517654 526255 519634 526280
rect 517132 526224 519634 526255
rect 519690 526224 519695 526280
rect 517132 526222 519695 526224
rect 517132 526195 517714 526222
rect 519629 526219 519695 526222
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 69013 517442 69079 517445
rect 71454 517442 72036 517455
rect 69013 517440 72036 517442
rect 69013 517384 69018 517440
rect 69074 517395 72036 517440
rect 69074 517384 71514 517395
rect 69013 517382 71514 517384
rect 69013 517379 69079 517382
rect 517132 515130 517714 515142
rect 519721 515130 519787 515133
rect 517132 515128 519787 515130
rect 517132 515082 519726 515128
rect 517654 515072 519726 515082
rect 519782 515072 519787 515128
rect 517654 515070 519787 515072
rect 519721 515067 519787 515070
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 69013 506562 69079 506565
rect 69013 506560 71514 506562
rect 69013 506504 69018 506560
rect 69074 506557 71514 506560
rect 69074 506504 72036 506557
rect 69013 506502 72036 506504
rect 69013 506499 69079 506502
rect 71454 506497 72036 506502
rect 519813 504114 519879 504117
rect 517654 504112 519879 504114
rect 517654 504056 519818 504112
rect 519874 504056 519879 504112
rect 517654 504054 519879 504056
rect 517654 504048 517714 504054
rect 519813 504051 519879 504054
rect 517132 503988 517714 504048
rect -960 501802 480 501892
rect 3601 501802 3667 501805
rect -960 501800 3667 501802
rect -960 501744 3606 501800
rect 3662 501744 3667 501800
rect -960 501742 3667 501744
rect -960 501652 480 501742
rect 3601 501739 3667 501742
rect 580165 497994 580231 497997
rect 583520 497994 584960 498084
rect 580165 497992 584960 497994
rect 580165 497936 580170 497992
rect 580226 497936 584960 497992
rect 580165 497934 584960 497936
rect 580165 497931 580231 497934
rect 583520 497844 584960 497934
rect 69013 495682 69079 495685
rect 69013 495680 71514 495682
rect 69013 495624 69018 495680
rect 69074 495660 71514 495680
rect 69074 495624 72036 495660
rect 69013 495622 72036 495624
rect 69013 495619 69079 495622
rect 71454 495600 72036 495622
rect 517132 492895 517714 492955
rect 517654 492826 517714 492895
rect 519537 492826 519603 492829
rect 517654 492824 519603 492826
rect 517654 492768 519542 492824
rect 519598 492768 519603 492824
rect 517654 492766 519603 492768
rect 519537 492763 519603 492766
rect -960 488746 480 488836
rect 3417 488746 3483 488749
rect -960 488744 3483 488746
rect -960 488688 3422 488744
rect 3478 488688 3483 488744
rect -960 488686 3483 488688
rect -960 488596 480 488686
rect 3417 488683 3483 488686
rect 69013 484802 69079 484805
rect 69013 484800 71514 484802
rect 69013 484744 69018 484800
rect 69074 484782 71514 484800
rect 69074 484744 72036 484782
rect 69013 484742 72036 484744
rect 69013 484739 69079 484742
rect 71454 484722 72036 484742
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 517132 481810 517714 481842
rect 519629 481810 519695 481813
rect 517132 481808 519695 481810
rect 517132 481782 519634 481808
rect 517654 481752 519634 481782
rect 519690 481752 519695 481808
rect 517654 481750 519695 481752
rect 519629 481747 519695 481750
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 69013 473922 69079 473925
rect 69013 473920 71514 473922
rect 69013 473864 69018 473920
rect 69074 473884 71514 473920
rect 69074 473864 72036 473884
rect 69013 473862 72036 473864
rect 69013 473859 69079 473862
rect 71454 473824 72036 473862
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 519721 470794 519787 470797
rect 517654 470792 519787 470794
rect 517654 470748 519726 470792
rect 517132 470736 519726 470748
rect 519782 470736 519787 470792
rect 517132 470734 519787 470736
rect 517132 470688 517714 470734
rect 519721 470731 519787 470734
rect 69013 463042 69079 463045
rect 69013 463040 71514 463042
rect 69013 462984 69018 463040
rect 69074 462986 71514 463040
rect 69074 462984 72036 462986
rect 69013 462982 72036 462984
rect 69013 462979 69079 462982
rect 71454 462926 72036 462982
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 519537 459642 519603 459645
rect 517654 459640 519603 459642
rect 517654 459635 519542 459640
rect 517132 459584 519542 459635
rect 519598 459584 519603 459640
rect 517132 459582 519603 459584
rect 517132 459575 517714 459582
rect 519537 459579 519603 459582
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 69013 452162 69079 452165
rect 69013 452160 71514 452162
rect 69013 452104 69018 452160
rect 69074 452108 71514 452160
rect 69074 452104 72036 452108
rect 69013 452102 72036 452104
rect 69013 452099 69079 452102
rect 71454 452048 72036 452102
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 519629 448626 519695 448629
rect 517654 448624 519695 448626
rect 517654 448568 519634 448624
rect 519690 448568 519695 448624
rect 517654 448566 519695 448568
rect 517654 448541 517714 448566
rect 519629 448563 519695 448566
rect 517132 448481 517714 448541
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 69013 441282 69079 441285
rect 69013 441280 71514 441282
rect 69013 441224 69018 441280
rect 69074 441224 71514 441280
rect 69013 441222 71514 441224
rect 69013 441219 69079 441222
rect 71454 441211 71514 441222
rect 71454 441151 72036 441211
rect 519537 437474 519603 437477
rect 517654 437472 519603 437474
rect 517654 437448 519542 437472
rect 517132 437416 519542 437448
rect 519598 437416 519603 437472
rect 517132 437414 519603 437416
rect 517132 437388 517714 437414
rect 519537 437411 519603 437414
rect -960 436658 480 436748
rect 3509 436658 3575 436661
rect -960 436656 3575 436658
rect -960 436600 3514 436656
rect 3570 436600 3575 436656
rect -960 436598 3575 436600
rect -960 436508 480 436598
rect 3509 436595 3575 436598
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 69013 430402 69079 430405
rect 69013 430400 71514 430402
rect 69013 430344 69018 430400
rect 69074 430344 71514 430400
rect 69013 430342 71514 430344
rect 69013 430339 69079 430342
rect 71454 430313 71514 430342
rect 71454 430253 72036 430313
rect 517132 426322 517714 426334
rect 519629 426322 519695 426325
rect 517132 426320 519695 426322
rect 517132 426274 519634 426320
rect 517654 426264 519634 426274
rect 519690 426264 519695 426320
rect 517654 426262 519695 426264
rect 519629 426259 519695 426262
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 69013 419386 69079 419389
rect 71454 419386 72036 419435
rect 69013 419384 72036 419386
rect 69013 419328 69018 419384
rect 69074 419375 72036 419384
rect 69074 419328 71514 419375
rect 69013 419326 71514 419328
rect 69013 419323 69079 419326
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 519537 415306 519603 415309
rect 517654 415304 519603 415306
rect 517654 415248 519542 415304
rect 519598 415248 519603 415304
rect 517654 415246 519603 415248
rect 517654 415241 517714 415246
rect 519537 415243 519603 415246
rect 517132 415181 517714 415241
rect -960 410546 480 410636
rect 3509 410546 3575 410549
rect -960 410544 3575 410546
rect -960 410488 3514 410544
rect 3570 410488 3575 410544
rect -960 410486 3575 410488
rect -960 410396 480 410486
rect 3509 410483 3575 410486
rect 69013 408642 69079 408645
rect 69013 408640 71514 408642
rect 69013 408584 69018 408640
rect 69074 408584 71514 408640
rect 69013 408582 71514 408584
rect 69013 408579 69079 408582
rect 71454 408538 71514 408582
rect 71454 408478 72036 408538
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 519629 404154 519695 404157
rect 517654 404152 519695 404154
rect 517654 404147 519634 404152
rect 517132 404096 519634 404147
rect 519690 404096 519695 404152
rect 517132 404094 519695 404096
rect 517132 404087 517714 404094
rect 519629 404091 519695 404094
rect 69013 397626 69079 397629
rect 71454 397626 72036 397640
rect 69013 397624 72036 397626
rect -960 397490 480 397580
rect 69013 397568 69018 397624
rect 69074 397580 72036 397624
rect 69074 397568 71514 397580
rect 69013 397566 71514 397568
rect 69013 397563 69079 397566
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 517132 393002 517714 393034
rect 519537 393002 519603 393005
rect 517132 393000 519603 393002
rect 517132 392974 519542 393000
rect 517654 392944 519542 392974
rect 519598 392944 519603 393000
rect 517654 392942 519603 392944
rect 519537 392939 519603 392942
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect 69013 386746 69079 386749
rect 71454 386746 72036 386762
rect 69013 386744 72036 386746
rect 69013 386688 69018 386744
rect 69074 386702 72036 386744
rect 69074 386688 71514 386702
rect 69013 386686 71514 386688
rect 69013 386683 69079 386686
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 519537 381986 519603 381989
rect 517654 381984 519603 381986
rect 517654 381940 519542 381984
rect 517132 381928 519542 381940
rect 519598 381928 519603 381984
rect 517132 381926 519603 381928
rect 517132 381880 517714 381926
rect 519537 381923 519603 381926
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 69013 375866 69079 375869
rect 69013 375864 71514 375866
rect 69013 375808 69018 375864
rect 69074 375808 72036 375864
rect 69013 375806 72036 375808
rect 69013 375803 69079 375806
rect 71454 375804 72036 375806
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 517132 370834 517714 370847
rect 519537 370834 519603 370837
rect 517132 370832 519603 370834
rect 517132 370787 519542 370832
rect 517654 370776 519542 370787
rect 519598 370776 519603 370832
rect 517654 370774 519603 370776
rect 519537 370771 519603 370774
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 69013 364986 69079 364989
rect 69013 364984 71514 364986
rect 69013 364928 69018 364984
rect 69074 364967 71514 364984
rect 583520 364972 584960 365062
rect 69074 364928 72036 364967
rect 69013 364926 72036 364928
rect 69013 364923 69079 364926
rect 71454 364907 72036 364926
rect 519353 359818 519419 359821
rect 517654 359816 519419 359818
rect 517654 359760 519358 359816
rect 519414 359760 519419 359816
rect 517654 359758 519419 359760
rect 517654 359734 517714 359758
rect 519353 359755 519419 359758
rect 517132 359674 517714 359734
rect -960 358458 480 358548
rect 3417 358458 3483 358461
rect -960 358456 3483 358458
rect -960 358400 3422 358456
rect 3478 358400 3483 358456
rect -960 358398 3483 358400
rect -960 358308 480 358398
rect 3417 358395 3483 358398
rect 69013 354106 69079 354109
rect 69013 354104 71514 354106
rect 69013 354048 69018 354104
rect 69074 354089 71514 354104
rect 69074 354048 72036 354089
rect 69013 354046 72036 354048
rect 69013 354043 69079 354046
rect 71454 354029 72036 354046
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 519813 348666 519879 348669
rect 517654 348664 519879 348666
rect 517654 348640 519818 348664
rect 517132 348608 519818 348640
rect 519874 348608 519879 348664
rect 517132 348606 519879 348608
rect 517132 348580 517714 348606
rect 519813 348603 519879 348606
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 69013 343226 69079 343229
rect 69013 343224 71514 343226
rect 69013 343168 69018 343224
rect 69074 343191 71514 343224
rect 69074 343168 72036 343191
rect 69013 343166 72036 343168
rect 69013 343163 69079 343166
rect 71454 343131 72036 343166
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 580165 338600 584960 338602
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect 517132 337514 517714 337546
rect 519997 337514 520063 337517
rect 517132 337512 520063 337514
rect 517132 337486 520002 337512
rect 517654 337456 520002 337486
rect 520058 337456 520063 337512
rect 517654 337454 520063 337456
rect 519997 337451 520063 337454
rect -960 332346 480 332436
rect 3417 332346 3483 332349
rect -960 332344 3483 332346
rect -960 332288 3422 332344
rect 3478 332288 3483 332344
rect -960 332286 3483 332288
rect -960 332196 480 332286
rect 3417 332283 3483 332286
rect 71454 332234 72036 332294
rect 69013 332210 69079 332213
rect 71454 332210 71514 332234
rect 69013 332208 71514 332210
rect 69013 332152 69018 332208
rect 69074 332152 71514 332208
rect 69013 332150 71514 332152
rect 69013 332147 69079 332150
rect 517132 326373 517714 326433
rect 517654 326362 517714 326373
rect 519353 326362 519419 326365
rect 517654 326360 519419 326362
rect 517654 326304 519358 326360
rect 519414 326304 519419 326360
rect 517654 326302 519419 326304
rect 519353 326299 519419 326302
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 71454 321356 72036 321416
rect 69013 321330 69079 321333
rect 71454 321330 71514 321356
rect 69013 321328 71514 321330
rect 69013 321272 69018 321328
rect 69074 321272 71514 321328
rect 69013 321270 71514 321272
rect 69013 321267 69079 321270
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 520181 315346 520247 315349
rect 517654 315344 520247 315346
rect 517654 315340 520186 315344
rect 517132 315288 520186 315340
rect 520242 315288 520247 315344
rect 517132 315286 520247 315288
rect 517132 315280 517714 315286
rect 520181 315283 520247 315286
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 71454 310458 72036 310518
rect 69013 310450 69079 310453
rect 71454 310450 71514 310458
rect 69013 310448 71514 310450
rect 69013 310392 69018 310448
rect 69074 310392 71514 310448
rect 69013 310390 71514 310392
rect 69013 310387 69079 310390
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 517132 304194 517714 304226
rect 519353 304194 519419 304197
rect 517132 304192 519419 304194
rect 517132 304166 519358 304192
rect 517654 304136 519358 304166
rect 519414 304136 519419 304192
rect 517654 304134 519419 304136
rect 519353 304131 519419 304134
rect 69013 299570 69079 299573
rect 71454 299570 72036 299620
rect 69013 299568 72036 299570
rect 69013 299512 69018 299568
rect 69074 299560 72036 299568
rect 69074 299512 71514 299560
rect 69013 299510 71514 299512
rect 69013 299507 69079 299510
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect 519537 293178 519603 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect 517654 293176 519603 293178
rect 517654 293133 519542 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 517132 293120 519542 293133
rect 519598 293120 519603 293176
rect 517132 293118 519603 293120
rect 517132 293073 517714 293118
rect 519537 293115 519603 293118
rect 69013 288690 69079 288693
rect 71454 288690 72036 288742
rect 69013 288688 72036 288690
rect 69013 288632 69018 288688
rect 69074 288682 72036 288688
rect 69074 288632 71514 288682
rect 69013 288630 71514 288632
rect 69013 288627 69079 288630
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 517132 282026 517714 282039
rect 519537 282026 519603 282029
rect 517132 282024 519603 282026
rect 517132 281979 519542 282024
rect 517654 281968 519542 281979
rect 519598 281968 519603 282024
rect 517654 281966 519603 281968
rect 519537 281963 519603 281966
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 69013 277810 69079 277813
rect 71454 277810 72036 277845
rect 69013 277808 72036 277810
rect 69013 277752 69018 277808
rect 69074 277785 72036 277808
rect 69074 277752 71514 277785
rect 69013 277750 71514 277752
rect 69013 277747 69079 277750
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 517132 270874 517714 270926
rect 519537 270874 519603 270877
rect 517132 270872 519603 270874
rect 517132 270866 519542 270872
rect 517654 270816 519542 270866
rect 519598 270816 519603 270872
rect 517654 270814 519603 270816
rect 519537 270811 519603 270814
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 69013 266930 69079 266933
rect 71454 266930 72036 266947
rect 69013 266928 72036 266930
rect 69013 266872 69018 266928
rect 69074 266887 72036 266928
rect 69074 266872 71514 266887
rect 69013 266870 71514 266872
rect 69013 266867 69079 266870
rect 519629 259858 519695 259861
rect 517654 259856 519695 259858
rect 517654 259832 519634 259856
rect 517132 259800 519634 259832
rect 519690 259800 519695 259856
rect 517132 259798 519695 259800
rect 517132 259772 517714 259798
rect 519629 259795 519695 259798
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 69013 256050 69079 256053
rect 71454 256050 72036 256069
rect 69013 256048 72036 256050
rect 69013 255992 69018 256048
rect 69074 256009 72036 256048
rect 69074 255992 71514 256009
rect 69013 255990 71514 255992
rect 69013 255987 69079 255990
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 517132 248706 517714 248739
rect 519537 248706 519603 248709
rect 517132 248704 519603 248706
rect 517132 248679 519542 248704
rect 517654 248648 519542 248679
rect 519598 248648 519603 248704
rect 517654 248646 519603 248648
rect 519537 248643 519603 248646
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 69013 245170 69079 245173
rect 71454 245170 72036 245172
rect 69013 245168 72036 245170
rect 69013 245112 69018 245168
rect 69074 245112 72036 245168
rect 69013 245110 71514 245112
rect 69013 245107 69079 245110
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 517132 237566 517714 237626
rect 517654 237554 517714 237566
rect 519629 237554 519695 237557
rect 517654 237552 519695 237554
rect 517654 237496 519634 237552
rect 519690 237496 519695 237552
rect 517654 237494 519695 237496
rect 519629 237491 519695 237494
rect 69013 234290 69079 234293
rect 69013 234288 71514 234290
rect 69013 234232 69018 234288
rect 69074 234274 71514 234288
rect 69074 234232 72036 234274
rect 69013 234230 72036 234232
rect 69013 234227 69079 234230
rect 71454 234214 72036 234230
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 519537 226538 519603 226541
rect 517654 226536 519603 226538
rect 517654 226532 519542 226536
rect 517132 226480 519542 226532
rect 519598 226480 519603 226536
rect 517132 226478 519603 226480
rect 517132 226472 517714 226478
rect 519537 226475 519603 226478
rect 69013 223410 69079 223413
rect 69013 223408 71514 223410
rect 69013 223352 69018 223408
rect 69074 223396 71514 223408
rect 69074 223352 72036 223396
rect 69013 223350 72036 223352
rect 69013 223347 69079 223350
rect 71454 223336 72036 223350
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 517132 215386 517714 215438
rect 519721 215386 519787 215389
rect 517132 215384 519787 215386
rect 517132 215378 519726 215384
rect 517654 215328 519726 215378
rect 519782 215328 519787 215384
rect 517654 215326 519787 215328
rect 519721 215323 519787 215326
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 69013 212530 69079 212533
rect 69013 212528 71514 212530
rect 69013 212472 69018 212528
rect 69074 212498 71514 212528
rect 69074 212472 72036 212498
rect 69013 212470 72036 212472
rect 69013 212467 69079 212470
rect 71454 212438 72036 212470
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 519629 204370 519695 204373
rect 517654 204368 519695 204370
rect 517654 204325 519634 204368
rect 517132 204312 519634 204325
rect 519690 204312 519695 204368
rect 517132 204310 519695 204312
rect 517132 204265 517714 204310
rect 519629 204307 519695 204310
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 69013 201650 69079 201653
rect 69013 201648 71514 201650
rect 69013 201592 69018 201648
rect 69074 201601 71514 201648
rect 69074 201592 72036 201601
rect 69013 201590 72036 201592
rect 69013 201587 69079 201590
rect 71454 201541 72036 201590
rect 517132 193218 517346 193232
rect 519537 193218 519603 193221
rect 517132 193216 519603 193218
rect 517132 193172 519542 193216
rect 517286 193160 519542 193172
rect 519598 193160 519603 193216
rect 517286 193158 519603 193160
rect 519537 193155 519603 193158
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 71454 190663 72036 190723
rect 69013 190634 69079 190637
rect 71454 190634 71514 190663
rect 69013 190632 71514 190634
rect 69013 190576 69018 190632
rect 69074 190576 71514 190632
rect 69013 190574 71514 190576
rect 69013 190571 69079 190574
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 517132 182066 517714 182118
rect 519721 182066 519787 182069
rect 517132 182064 519787 182066
rect 517132 182058 519726 182064
rect 517654 182008 519726 182058
rect 519782 182008 519787 182064
rect 517654 182006 519787 182008
rect 519721 182003 519787 182006
rect 71454 179765 72036 179825
rect 69013 179754 69079 179757
rect 71454 179754 71514 179765
rect 69013 179752 71514 179754
rect 69013 179696 69018 179752
rect 69074 179696 71514 179752
rect 69013 179694 71514 179696
rect 69013 179691 69079 179694
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 3509 175946 3575 175949
rect -960 175944 3575 175946
rect -960 175888 3514 175944
rect 3570 175888 3575 175944
rect -960 175886 3575 175888
rect -960 175796 480 175886
rect 3509 175883 3575 175886
rect 519629 171050 519695 171053
rect 517654 171048 519695 171050
rect 517654 171025 519634 171048
rect 517132 170992 519634 171025
rect 519690 170992 519695 171048
rect 517132 170990 519695 170992
rect 517132 170965 517714 170990
rect 519629 170987 519695 170990
rect 69013 168874 69079 168877
rect 71454 168874 72036 168928
rect 69013 168872 72036 168874
rect 69013 168816 69018 168872
rect 69074 168868 72036 168872
rect 69074 168816 71514 168868
rect 69013 168814 71514 168816
rect 69013 168811 69079 168814
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 517132 159898 517714 159931
rect 519537 159898 519603 159901
rect 517132 159896 519603 159898
rect 517132 159871 519542 159896
rect 517654 159840 519542 159871
rect 519598 159840 519603 159896
rect 517654 159838 519603 159840
rect 519537 159835 519603 159838
rect 69013 157994 69079 157997
rect 71454 157994 72036 158050
rect 69013 157992 72036 157994
rect 69013 157936 69018 157992
rect 69074 157990 72036 157992
rect 69074 157936 71514 157990
rect 69013 157934 71514 157936
rect 69013 157931 69079 157934
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 517132 148758 517714 148818
rect 517654 148746 517714 148758
rect 519813 148746 519879 148749
rect 517654 148744 519879 148746
rect 517654 148688 519818 148744
rect 519874 148688 519879 148744
rect 517654 148686 519879 148688
rect 519813 148683 519879 148686
rect 69013 147114 69079 147117
rect 71454 147114 72036 147152
rect 69013 147112 72036 147114
rect 69013 147056 69018 147112
rect 69074 147092 72036 147112
rect 69074 147056 71514 147092
rect 69013 147054 71514 147056
rect 69013 147051 69079 147054
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 519721 137730 519787 137733
rect 517654 137728 519787 137730
rect 517654 137724 519726 137728
rect 517132 137672 519726 137724
rect 519782 137672 519787 137728
rect 517132 137670 519787 137672
rect 517132 137664 517714 137670
rect 519721 137667 519787 137670
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 69013 136234 69079 136237
rect 71454 136234 72036 136254
rect 69013 136232 72036 136234
rect 69013 136176 69018 136232
rect 69074 136194 72036 136232
rect 69074 136176 71514 136194
rect 69013 136174 71514 136176
rect 69013 136171 69079 136174
rect 517132 126578 517714 126631
rect 519629 126578 519695 126581
rect 517132 126576 519695 126578
rect 517132 126571 519634 126576
rect 517654 126520 519634 126571
rect 519690 126520 519695 126576
rect 517654 126518 519695 126520
rect 519629 126515 519695 126518
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 69013 125354 69079 125357
rect 71454 125354 72036 125376
rect 69013 125352 72036 125354
rect 69013 125296 69018 125352
rect 69074 125316 72036 125352
rect 69074 125296 71514 125316
rect 69013 125294 71514 125296
rect 69013 125291 69079 125294
rect -960 123722 480 123812
rect 3417 123722 3483 123725
rect -960 123720 3483 123722
rect -960 123664 3422 123720
rect 3478 123664 3483 123720
rect -960 123662 3483 123664
rect -960 123572 480 123662
rect 3417 123659 3483 123662
rect 519537 115562 519603 115565
rect 517654 115560 519603 115562
rect 517654 115518 519542 115560
rect 517132 115504 519542 115518
rect 519598 115504 519603 115560
rect 517132 115502 519603 115504
rect 517132 115458 517714 115502
rect 519537 115499 519603 115502
rect 69013 114474 69079 114477
rect 71454 114474 72036 114479
rect 69013 114472 72036 114474
rect 69013 114416 69018 114472
rect 69074 114419 72036 114472
rect 69074 114416 71514 114419
rect 69013 114414 71514 114416
rect 69013 114411 69079 114414
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3693 110666 3759 110669
rect -960 110664 3759 110666
rect -960 110608 3698 110664
rect 3754 110608 3759 110664
rect -960 110606 3759 110608
rect -960 110516 480 110606
rect 3693 110603 3759 110606
rect 517132 104410 517714 104424
rect 519905 104410 519971 104413
rect 517132 104408 519971 104410
rect 517132 104364 519910 104408
rect 517654 104352 519910 104364
rect 519966 104352 519971 104408
rect 517654 104350 519971 104352
rect 519905 104347 519971 104350
rect 69013 103594 69079 103597
rect 69013 103592 71514 103594
rect 69013 103536 69018 103592
rect 69074 103581 71514 103592
rect 69074 103536 72036 103581
rect 69013 103534 72036 103536
rect 69013 103531 69079 103534
rect 71454 103521 72036 103534
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 517132 93270 517714 93330
rect 517654 93258 517714 93270
rect 519813 93258 519879 93261
rect 517654 93256 519879 93258
rect 517654 93200 519818 93256
rect 519874 93200 519879 93256
rect 517654 93198 519879 93200
rect 519813 93195 519879 93198
rect 69013 92714 69079 92717
rect 69013 92712 71514 92714
rect 69013 92656 69018 92712
rect 69074 92703 71514 92712
rect 69074 92656 72036 92703
rect 69013 92654 72036 92656
rect 69013 92651 69079 92654
rect 71454 92643 72036 92654
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 519721 82242 519787 82245
rect 517654 82240 519787 82242
rect 517654 82217 519726 82240
rect 517132 82184 519726 82217
rect 519782 82184 519787 82240
rect 517132 82182 519787 82184
rect 517132 82157 517714 82182
rect 519721 82179 519787 82182
rect 69013 81834 69079 81837
rect 69013 81832 71514 81834
rect 69013 81776 69018 81832
rect 69074 81806 71514 81832
rect 69074 81776 72036 81806
rect 69013 81774 72036 81776
rect 69013 81771 69079 81774
rect 71454 81746 72036 81774
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 517132 71090 517714 71124
rect 519629 71090 519695 71093
rect 517132 71088 519695 71090
rect 517132 71064 519634 71088
rect 517654 71032 519634 71064
rect 519690 71032 519695 71088
rect 517654 71030 519695 71032
rect 519629 71027 519695 71030
rect 71454 70848 72036 70908
rect 69013 70818 69079 70821
rect 71454 70818 71514 70848
rect 69013 70816 71514 70818
rect 69013 70760 69018 70816
rect 69074 70760 71514 70816
rect 69013 70758 71514 70760
rect 69013 70755 69079 70758
rect 517132 60482 517714 60520
rect 519537 60482 519603 60485
rect 517132 60480 519603 60482
rect 517132 60460 519542 60480
rect 517654 60424 519542 60460
rect 519598 60424 519603 60480
rect 517654 60422 519603 60424
rect 519537 60419 519603 60422
rect 71454 60225 72036 60285
rect 69013 60210 69079 60213
rect 71454 60210 71514 60225
rect 69013 60208 71514 60210
rect 69013 60152 69018 60208
rect 69074 60152 71514 60208
rect 69013 60150 71514 60152
rect 69013 60147 69079 60150
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3785 58578 3851 58581
rect -960 58576 3851 58578
rect -960 58520 3790 58576
rect 3846 58520 3851 58576
rect -960 58518 3851 58520
rect -960 58428 480 58518
rect 3785 58515 3851 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3601 32466 3667 32469
rect -960 32464 3667 32466
rect -960 32408 3606 32464
rect 3662 32408 3667 32464
rect -960 32406 3667 32408
rect -960 32316 480 32406
rect 3601 32403 3667 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 19425 3770 19491 3773
rect 133965 3770 134031 3773
rect 19425 3768 134031 3770
rect 19425 3712 19430 3768
rect 19486 3712 133970 3768
rect 134026 3712 134031 3768
rect 19425 3710 134031 3712
rect 19425 3707 19491 3710
rect 133965 3707 134031 3710
rect 362309 3770 362375 3773
rect 458265 3770 458331 3773
rect 362309 3768 458331 3770
rect 362309 3712 362314 3768
rect 362370 3712 458270 3768
rect 458326 3712 458331 3768
rect 362309 3710 458331 3712
rect 362309 3707 362375 3710
rect 458265 3707 458331 3710
rect 20621 3634 20687 3637
rect 162945 3634 163011 3637
rect 20621 3632 163011 3634
rect 20621 3576 20626 3632
rect 20682 3576 162950 3632
rect 163006 3576 163011 3632
rect 20621 3574 163011 3576
rect 20621 3571 20687 3574
rect 162945 3571 163011 3574
rect 358721 3634 358787 3637
rect 456793 3634 456859 3637
rect 358721 3632 456859 3634
rect 358721 3576 358726 3632
rect 358782 3576 456798 3632
rect 456854 3576 456859 3632
rect 358721 3574 456859 3576
rect 358721 3571 358787 3574
rect 456793 3571 456859 3574
rect 11145 3498 11211 3501
rect 161565 3498 161631 3501
rect 11145 3496 161631 3498
rect 11145 3440 11150 3496
rect 11206 3440 161570 3496
rect 161626 3440 161631 3496
rect 11145 3438 161631 3440
rect 11145 3435 11211 3438
rect 161565 3435 161631 3438
rect 355225 3498 355291 3501
rect 455597 3498 455663 3501
rect 355225 3496 455663 3498
rect 355225 3440 355230 3496
rect 355286 3440 455602 3496
rect 455658 3440 455663 3496
rect 355225 3438 455663 3440
rect 355225 3435 355291 3438
rect 455597 3435 455663 3438
rect 516041 3498 516107 3501
rect 580993 3498 581059 3501
rect 516041 3496 581059 3498
rect 516041 3440 516046 3496
rect 516102 3440 580998 3496
rect 581054 3440 581059 3496
rect 516041 3438 581059 3440
rect 516041 3435 516107 3438
rect 580993 3435 581059 3438
rect 5257 3362 5323 3365
rect 165705 3362 165771 3365
rect 5257 3360 165771 3362
rect 5257 3304 5262 3360
rect 5318 3304 165710 3360
rect 165766 3304 165771 3360
rect 5257 3302 165771 3304
rect 5257 3299 5323 3302
rect 165705 3299 165771 3302
rect 351637 3362 351703 3365
rect 455505 3362 455571 3365
rect 351637 3360 455571 3362
rect 351637 3304 351642 3360
rect 351698 3304 455510 3360
rect 455566 3304 455571 3360
rect 351637 3302 455571 3304
rect 351637 3299 351703 3302
rect 455505 3299 455571 3302
rect 517421 3362 517487 3365
rect 583385 3362 583451 3365
rect 517421 3360 583451 3362
rect 517421 3304 517426 3360
rect 517482 3304 583390 3360
rect 583446 3304 583451 3360
rect 517421 3302 583451 3304
rect 517421 3299 517487 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 641020 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 641020 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 641020 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 641020 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 641020 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 641020 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 641020 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 641020 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 641020 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 641020 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 641020 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 641020 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 641020 128414 668898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 641020 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 641020 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 641020 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 641020 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 641020 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 641020 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 641020 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 641020 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 641020 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 641020 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 641020 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 641020 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 641020 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 641020 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 641020 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 641020 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 641020 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 641020 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 641020 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 641020 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 641020 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 641020 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 641020 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 641020 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 641020 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 641020 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 641020 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 641020 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 641020 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 641020 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 641020 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 641020 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 641020 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 641020 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 641020 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 641020 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 641020 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 641020 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 641020 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 641020 308414 668898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 641020 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 641020 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 641020 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 641020 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 641020 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 641020 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 641020 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 641020 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 641020 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 641020 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 641020 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 641020 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 641020 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 641020 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 641020 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 641020 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 641020 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 641020 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 641020 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 641020 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 641020 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 641020 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 641020 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 641020 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 641020 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 641020 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 641020 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 641020 434414 650898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 641020 438134 654618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 641020 441854 658338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 641020 445574 662058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 641020 452414 668898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 641020 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 641020 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 641020 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 641020 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 641020 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 641020 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 641020 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 641020 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 641020 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 641020 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 641020 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 641020 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 641020 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 641020 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 641020 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 289457 615454 289857 615486
rect 289457 615218 289539 615454
rect 289775 615218 289857 615454
rect 289457 615134 289857 615218
rect 289457 614898 289539 615134
rect 289775 614898 289857 615134
rect 289457 614866 289857 614898
rect 505845 615454 506245 615486
rect 505845 615218 505927 615454
rect 506163 615218 506245 615454
rect 505845 615134 506245 615218
rect 505845 614898 505927 615134
rect 506163 614898 506245 615134
rect 505845 614866 506245 614898
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 288697 597454 289097 597486
rect 288697 597218 288779 597454
rect 289015 597218 289097 597454
rect 288697 597134 289097 597218
rect 288697 596898 288779 597134
rect 289015 596898 289097 597134
rect 288697 596866 289097 596898
rect 293911 597454 294259 597486
rect 293911 597218 293967 597454
rect 294203 597218 294259 597454
rect 293911 597134 294259 597218
rect 293911 596898 293967 597134
rect 294203 596898 294259 597134
rect 293911 596866 294259 596898
rect 388975 597454 389323 597486
rect 388975 597218 389031 597454
rect 389267 597218 389323 597454
rect 388975 597134 389323 597218
rect 388975 596898 389031 597134
rect 389267 596898 389323 597134
rect 388975 596866 389323 596898
rect 406339 597454 406687 597486
rect 406339 597218 406395 597454
rect 406631 597218 406687 597454
rect 406339 597134 406687 597218
rect 406339 596898 406395 597134
rect 406631 596898 406687 597134
rect 406339 596866 406687 596898
rect 501403 597454 501751 597486
rect 501403 597218 501459 597454
rect 501695 597218 501751 597454
rect 501403 597134 501751 597218
rect 501403 596898 501459 597134
rect 501695 596898 501751 597134
rect 501403 596866 501751 596898
rect 506605 597454 507005 597486
rect 506605 597218 506687 597454
rect 506923 597218 507005 597454
rect 506605 597134 507005 597218
rect 506605 596898 506687 597134
rect 506923 596898 507005 597134
rect 506605 596866 507005 596898
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 289457 579454 289857 579486
rect 289457 579218 289539 579454
rect 289775 579218 289857 579454
rect 289457 579134 289857 579218
rect 289457 578898 289539 579134
rect 289775 578898 289857 579134
rect 289457 578866 289857 578898
rect 294591 579454 294939 579486
rect 294591 579218 294647 579454
rect 294883 579218 294939 579454
rect 294591 579134 294939 579218
rect 294591 578898 294647 579134
rect 294883 578898 294939 579134
rect 294591 578866 294939 578898
rect 388295 579454 388643 579486
rect 388295 579218 388351 579454
rect 388587 579218 388643 579454
rect 388295 579134 388643 579218
rect 388295 578898 388351 579134
rect 388587 578898 388643 579134
rect 388295 578866 388643 578898
rect 407019 579454 407367 579486
rect 407019 579218 407075 579454
rect 407311 579218 407367 579454
rect 407019 579134 407367 579218
rect 407019 578898 407075 579134
rect 407311 578898 407367 579134
rect 407019 578866 407367 578898
rect 500723 579454 501071 579486
rect 500723 579218 500779 579454
rect 501015 579218 501071 579454
rect 500723 579134 501071 579218
rect 500723 578898 500779 579134
rect 501015 578898 501071 579134
rect 500723 578866 501071 578898
rect 505845 579454 506245 579486
rect 505845 579218 505927 579454
rect 506163 579218 506245 579454
rect 505845 579134 506245 579218
rect 505845 578898 505927 579134
rect 506163 578898 506245 579134
rect 505845 578866 506245 578898
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 288697 561454 289097 561486
rect 288697 561218 288779 561454
rect 289015 561218 289097 561454
rect 288697 561134 289097 561218
rect 288697 560898 288779 561134
rect 289015 560898 289097 561134
rect 288697 560866 289097 560898
rect 293911 561454 294259 561486
rect 293911 561218 293967 561454
rect 294203 561218 294259 561454
rect 293911 561134 294259 561218
rect 293911 560898 293967 561134
rect 294203 560898 294259 561134
rect 293911 560866 294259 560898
rect 388975 561454 389323 561486
rect 388975 561218 389031 561454
rect 389267 561218 389323 561454
rect 388975 561134 389323 561218
rect 388975 560898 389031 561134
rect 389267 560898 389323 561134
rect 388975 560866 389323 560898
rect 406339 561454 406687 561486
rect 406339 561218 406395 561454
rect 406631 561218 406687 561454
rect 406339 561134 406687 561218
rect 406339 560898 406395 561134
rect 406631 560898 406687 561134
rect 406339 560866 406687 560898
rect 501403 561454 501751 561486
rect 501403 561218 501459 561454
rect 501695 561218 501751 561454
rect 501403 561134 501751 561218
rect 501403 560898 501459 561134
rect 501695 560898 501751 561134
rect 501403 560866 501751 560898
rect 506605 561454 507005 561486
rect 506605 561218 506687 561454
rect 506923 561218 507005 561454
rect 506605 561134 507005 561218
rect 506605 560898 506687 561134
rect 506923 560898 507005 561134
rect 506605 560866 507005 560898
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 289457 543454 289857 543486
rect 289457 543218 289539 543454
rect 289775 543218 289857 543454
rect 289457 543134 289857 543218
rect 289457 542898 289539 543134
rect 289775 542898 289857 543134
rect 289457 542866 289857 542898
rect 294591 543454 294939 543486
rect 294591 543218 294647 543454
rect 294883 543218 294939 543454
rect 294591 543134 294939 543218
rect 294591 542898 294647 543134
rect 294883 542898 294939 543134
rect 294591 542866 294939 542898
rect 388295 543454 388643 543486
rect 388295 543218 388351 543454
rect 388587 543218 388643 543454
rect 388295 543134 388643 543218
rect 388295 542898 388351 543134
rect 388587 542898 388643 543134
rect 388295 542866 388643 542898
rect 407019 543454 407367 543486
rect 407019 543218 407075 543454
rect 407311 543218 407367 543454
rect 407019 543134 407367 543218
rect 407019 542898 407075 543134
rect 407311 542898 407367 543134
rect 407019 542866 407367 542898
rect 500723 543454 501071 543486
rect 500723 543218 500779 543454
rect 501015 543218 501071 543454
rect 500723 543134 501071 543218
rect 500723 542898 500779 543134
rect 501015 542898 501071 543134
rect 500723 542866 501071 542898
rect 505845 543454 506245 543486
rect 505845 543218 505927 543454
rect 506163 543218 506245 543454
rect 505845 543134 506245 543218
rect 505845 542898 505927 543134
rect 506163 542898 506245 543134
rect 505845 542866 506245 542898
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 288213 489454 288561 489486
rect 288213 489218 288269 489454
rect 288505 489218 288561 489454
rect 288213 489134 288561 489218
rect 288213 488898 288269 489134
rect 288505 488898 288561 489134
rect 288213 488866 288561 488898
rect 383277 489454 383625 489486
rect 383277 489218 383333 489454
rect 383569 489218 383625 489454
rect 383277 489134 383625 489218
rect 383277 488898 383333 489134
rect 383569 488898 383625 489134
rect 383277 488866 383625 488898
rect 412183 489454 412531 489486
rect 412183 489218 412239 489454
rect 412475 489218 412531 489454
rect 412183 489134 412531 489218
rect 412183 488898 412239 489134
rect 412475 488898 412531 489134
rect 412183 488866 412531 488898
rect 507247 489454 507595 489486
rect 507247 489218 507303 489454
rect 507539 489218 507595 489454
rect 507247 489134 507595 489218
rect 507247 488898 507303 489134
rect 507539 488898 507595 489134
rect 507247 488866 507595 488898
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 288893 471454 289241 471486
rect 288893 471218 288949 471454
rect 289185 471218 289241 471454
rect 288893 471134 289241 471218
rect 288893 470898 288949 471134
rect 289185 470898 289241 471134
rect 288893 470866 289241 470898
rect 382597 471454 382945 471486
rect 382597 471218 382653 471454
rect 382889 471218 382945 471454
rect 382597 471134 382945 471218
rect 382597 470898 382653 471134
rect 382889 470898 382945 471134
rect 382597 470866 382945 470898
rect 412863 471454 413211 471486
rect 412863 471218 412919 471454
rect 413155 471218 413211 471454
rect 412863 471134 413211 471218
rect 412863 470898 412919 471134
rect 413155 470898 413211 471134
rect 412863 470866 413211 470898
rect 506567 471454 506915 471486
rect 506567 471218 506623 471454
rect 506859 471218 506915 471454
rect 506567 471134 506915 471218
rect 506567 470898 506623 471134
rect 506859 470898 506915 471134
rect 506567 470866 506915 470898
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 288213 453454 288561 453486
rect 288213 453218 288269 453454
rect 288505 453218 288561 453454
rect 288213 453134 288561 453218
rect 288213 452898 288269 453134
rect 288505 452898 288561 453134
rect 288213 452866 288561 452898
rect 383277 453454 383625 453486
rect 383277 453218 383333 453454
rect 383569 453218 383625 453454
rect 383277 453134 383625 453218
rect 383277 452898 383333 453134
rect 383569 452898 383625 453134
rect 383277 452866 383625 452898
rect 412183 453454 412531 453486
rect 412183 453218 412239 453454
rect 412475 453218 412531 453454
rect 412183 453134 412531 453218
rect 412183 452898 412239 453134
rect 412475 452898 412531 453134
rect 412183 452866 412531 452898
rect 507247 453454 507595 453486
rect 507247 453218 507303 453454
rect 507539 453218 507595 453454
rect 507247 453134 507595 453218
rect 507247 452898 507303 453134
rect 507539 452898 507595 453134
rect 507247 452866 507595 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 288893 435454 289241 435486
rect 288893 435218 288949 435454
rect 289185 435218 289241 435454
rect 288893 435134 289241 435218
rect 288893 434898 288949 435134
rect 289185 434898 289241 435134
rect 288893 434866 289241 434898
rect 382597 435454 382945 435486
rect 382597 435218 382653 435454
rect 382889 435218 382945 435454
rect 382597 435134 382945 435218
rect 382597 434898 382653 435134
rect 382889 434898 382945 435134
rect 382597 434866 382945 434898
rect 412863 435454 413211 435486
rect 412863 435218 412919 435454
rect 413155 435218 413211 435454
rect 412863 435134 413211 435218
rect 412863 434898 412919 435134
rect 413155 434898 413211 435134
rect 412863 434866 413211 434898
rect 506567 435454 506915 435486
rect 506567 435218 506623 435454
rect 506859 435218 506915 435454
rect 506567 435134 506915 435218
rect 506567 434898 506623 435134
rect 506859 434898 506915 435134
rect 506567 434866 506915 434898
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 288893 399454 289241 399486
rect 288893 399218 288949 399454
rect 289185 399218 289241 399454
rect 288893 399134 289241 399218
rect 288893 398898 288949 399134
rect 289185 398898 289241 399134
rect 288893 398866 289241 398898
rect 382597 399454 382945 399486
rect 382597 399218 382653 399454
rect 382889 399218 382945 399454
rect 382597 399134 382945 399218
rect 382597 398898 382653 399134
rect 382889 398898 382945 399134
rect 382597 398866 382945 398898
rect 412863 399454 413211 399486
rect 412863 399218 412919 399454
rect 413155 399218 413211 399454
rect 412863 399134 413211 399218
rect 412863 398898 412919 399134
rect 413155 398898 413211 399134
rect 412863 398866 413211 398898
rect 506567 399454 506915 399486
rect 506567 399218 506623 399454
rect 506859 399218 506915 399454
rect 506567 399134 506915 399218
rect 506567 398898 506623 399134
rect 506859 398898 506915 399134
rect 506567 398866 506915 398898
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 288213 381454 288561 381486
rect 288213 381218 288269 381454
rect 288505 381218 288561 381454
rect 288213 381134 288561 381218
rect 288213 380898 288269 381134
rect 288505 380898 288561 381134
rect 288213 380866 288561 380898
rect 383277 381454 383625 381486
rect 383277 381218 383333 381454
rect 383569 381218 383625 381454
rect 383277 381134 383625 381218
rect 383277 380898 383333 381134
rect 383569 380898 383625 381134
rect 383277 380866 383625 380898
rect 412183 381454 412531 381486
rect 412183 381218 412239 381454
rect 412475 381218 412531 381454
rect 412183 381134 412531 381218
rect 412183 380898 412239 381134
rect 412475 380898 412531 381134
rect 412183 380866 412531 380898
rect 507247 381454 507595 381486
rect 507247 381218 507303 381454
rect 507539 381218 507595 381454
rect 507247 381134 507595 381218
rect 507247 380898 507303 381134
rect 507539 380898 507595 381134
rect 507247 380866 507595 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 288893 363454 289241 363486
rect 288893 363218 288949 363454
rect 289185 363218 289241 363454
rect 288893 363134 289241 363218
rect 288893 362898 288949 363134
rect 289185 362898 289241 363134
rect 288893 362866 289241 362898
rect 382597 363454 382945 363486
rect 382597 363218 382653 363454
rect 382889 363218 382945 363454
rect 382597 363134 382945 363218
rect 382597 362898 382653 363134
rect 382889 362898 382945 363134
rect 382597 362866 382945 362898
rect 412863 363454 413211 363486
rect 412863 363218 412919 363454
rect 413155 363218 413211 363454
rect 412863 363134 413211 363218
rect 412863 362898 412919 363134
rect 413155 362898 413211 363134
rect 412863 362866 413211 362898
rect 506567 363454 506915 363486
rect 506567 363218 506623 363454
rect 506859 363218 506915 363454
rect 506567 363134 506915 363218
rect 506567 362898 506623 363134
rect 506859 362898 506915 363134
rect 506567 362866 506915 362898
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 288213 345454 288561 345486
rect 288213 345218 288269 345454
rect 288505 345218 288561 345454
rect 288213 345134 288561 345218
rect 288213 344898 288269 345134
rect 288505 344898 288561 345134
rect 288213 344866 288561 344898
rect 383277 345454 383625 345486
rect 383277 345218 383333 345454
rect 383569 345218 383625 345454
rect 383277 345134 383625 345218
rect 383277 344898 383333 345134
rect 383569 344898 383625 345134
rect 383277 344866 383625 344898
rect 412183 345454 412531 345486
rect 412183 345218 412239 345454
rect 412475 345218 412531 345454
rect 412183 345134 412531 345218
rect 412183 344898 412239 345134
rect 412475 344898 412531 345134
rect 412183 344866 412531 344898
rect 507247 345454 507595 345486
rect 507247 345218 507303 345454
rect 507539 345218 507595 345454
rect 507247 345134 507595 345218
rect 507247 344898 507303 345134
rect 507539 344898 507595 345134
rect 507247 344866 507595 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 288893 291454 289241 291486
rect 288893 291218 288949 291454
rect 289185 291218 289241 291454
rect 288893 291134 289241 291218
rect 288893 290898 288949 291134
rect 289185 290898 289241 291134
rect 288893 290866 289241 290898
rect 382597 291454 382945 291486
rect 382597 291218 382653 291454
rect 382889 291218 382945 291454
rect 382597 291134 382945 291218
rect 382597 290898 382653 291134
rect 382889 290898 382945 291134
rect 382597 290866 382945 290898
rect 412863 291454 413211 291486
rect 412863 291218 412919 291454
rect 413155 291218 413211 291454
rect 412863 291134 413211 291218
rect 412863 290898 412919 291134
rect 413155 290898 413211 291134
rect 412863 290866 413211 290898
rect 506567 291454 506915 291486
rect 506567 291218 506623 291454
rect 506859 291218 506915 291454
rect 506567 291134 506915 291218
rect 506567 290898 506623 291134
rect 506859 290898 506915 291134
rect 506567 290866 506915 290898
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 288213 273454 288561 273486
rect 288213 273218 288269 273454
rect 288505 273218 288561 273454
rect 288213 273134 288561 273218
rect 288213 272898 288269 273134
rect 288505 272898 288561 273134
rect 288213 272866 288561 272898
rect 383277 273454 383625 273486
rect 383277 273218 383333 273454
rect 383569 273218 383625 273454
rect 383277 273134 383625 273218
rect 383277 272898 383333 273134
rect 383569 272898 383625 273134
rect 383277 272866 383625 272898
rect 412183 273454 412531 273486
rect 412183 273218 412239 273454
rect 412475 273218 412531 273454
rect 412183 273134 412531 273218
rect 412183 272898 412239 273134
rect 412475 272898 412531 273134
rect 412183 272866 412531 272898
rect 507247 273454 507595 273486
rect 507247 273218 507303 273454
rect 507539 273218 507595 273454
rect 507247 273134 507595 273218
rect 507247 272898 507303 273134
rect 507539 272898 507595 273134
rect 507247 272866 507595 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 288893 255454 289241 255486
rect 288893 255218 288949 255454
rect 289185 255218 289241 255454
rect 288893 255134 289241 255218
rect 288893 254898 288949 255134
rect 289185 254898 289241 255134
rect 288893 254866 289241 254898
rect 382597 255454 382945 255486
rect 382597 255218 382653 255454
rect 382889 255218 382945 255454
rect 382597 255134 382945 255218
rect 382597 254898 382653 255134
rect 382889 254898 382945 255134
rect 382597 254866 382945 254898
rect 412863 255454 413211 255486
rect 412863 255218 412919 255454
rect 413155 255218 413211 255454
rect 412863 255134 413211 255218
rect 412863 254898 412919 255134
rect 413155 254898 413211 255134
rect 412863 254866 413211 254898
rect 506567 255454 506915 255486
rect 506567 255218 506623 255454
rect 506859 255218 506915 255454
rect 506567 255134 506915 255218
rect 506567 254898 506623 255134
rect 506859 254898 506915 255134
rect 506567 254866 506915 254898
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 288213 237454 288561 237486
rect 288213 237218 288269 237454
rect 288505 237218 288561 237454
rect 288213 237134 288561 237218
rect 288213 236898 288269 237134
rect 288505 236898 288561 237134
rect 288213 236866 288561 236898
rect 383277 237454 383625 237486
rect 383277 237218 383333 237454
rect 383569 237218 383625 237454
rect 383277 237134 383625 237218
rect 383277 236898 383333 237134
rect 383569 236898 383625 237134
rect 383277 236866 383625 236898
rect 412183 237454 412531 237486
rect 412183 237218 412239 237454
rect 412475 237218 412531 237454
rect 412183 237134 412531 237218
rect 412183 236898 412239 237134
rect 412475 236898 412531 237134
rect 412183 236866 412531 236898
rect 507247 237454 507595 237486
rect 507247 237218 507303 237454
rect 507539 237218 507595 237454
rect 507247 237134 507595 237218
rect 507247 236898 507303 237134
rect 507539 236898 507595 237134
rect 507247 236866 507595 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 288213 201454 288561 201486
rect 288213 201218 288269 201454
rect 288505 201218 288561 201454
rect 288213 201134 288561 201218
rect 288213 200898 288269 201134
rect 288505 200898 288561 201134
rect 288213 200866 288561 200898
rect 383277 201454 383625 201486
rect 383277 201218 383333 201454
rect 383569 201218 383625 201454
rect 383277 201134 383625 201218
rect 383277 200898 383333 201134
rect 383569 200898 383625 201134
rect 383277 200866 383625 200898
rect 412183 201454 412531 201486
rect 412183 201218 412239 201454
rect 412475 201218 412531 201454
rect 412183 201134 412531 201218
rect 412183 200898 412239 201134
rect 412475 200898 412531 201134
rect 412183 200866 412531 200898
rect 507247 201454 507595 201486
rect 507247 201218 507303 201454
rect 507539 201218 507595 201454
rect 507247 201134 507595 201218
rect 507247 200898 507303 201134
rect 507539 200898 507595 201134
rect 507247 200866 507595 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 288893 183454 289241 183486
rect 288893 183218 288949 183454
rect 289185 183218 289241 183454
rect 288893 183134 289241 183218
rect 288893 182898 288949 183134
rect 289185 182898 289241 183134
rect 288893 182866 289241 182898
rect 382597 183454 382945 183486
rect 382597 183218 382653 183454
rect 382889 183218 382945 183454
rect 382597 183134 382945 183218
rect 382597 182898 382653 183134
rect 382889 182898 382945 183134
rect 382597 182866 382945 182898
rect 412863 183454 413211 183486
rect 412863 183218 412919 183454
rect 413155 183218 413211 183454
rect 412863 183134 413211 183218
rect 412863 182898 412919 183134
rect 413155 182898 413211 183134
rect 412863 182866 413211 182898
rect 506567 183454 506915 183486
rect 506567 183218 506623 183454
rect 506859 183218 506915 183454
rect 506567 183134 506915 183218
rect 506567 182898 506623 183134
rect 506859 182898 506915 183134
rect 506567 182866 506915 182898
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 288213 165454 288561 165486
rect 288213 165218 288269 165454
rect 288505 165218 288561 165454
rect 288213 165134 288561 165218
rect 288213 164898 288269 165134
rect 288505 164898 288561 165134
rect 288213 164866 288561 164898
rect 383277 165454 383625 165486
rect 383277 165218 383333 165454
rect 383569 165218 383625 165454
rect 383277 165134 383625 165218
rect 383277 164898 383333 165134
rect 383569 164898 383625 165134
rect 383277 164866 383625 164898
rect 412183 165454 412531 165486
rect 412183 165218 412239 165454
rect 412475 165218 412531 165454
rect 412183 165134 412531 165218
rect 412183 164898 412239 165134
rect 412475 164898 412531 165134
rect 412183 164866 412531 164898
rect 507247 165454 507595 165486
rect 507247 165218 507303 165454
rect 507539 165218 507595 165454
rect 507247 165134 507595 165218
rect 507247 164898 507303 165134
rect 507539 164898 507595 165134
rect 507247 164866 507595 164898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 288893 147454 289241 147486
rect 288893 147218 288949 147454
rect 289185 147218 289241 147454
rect 288893 147134 289241 147218
rect 288893 146898 288949 147134
rect 289185 146898 289241 147134
rect 288893 146866 289241 146898
rect 382597 147454 382945 147486
rect 382597 147218 382653 147454
rect 382889 147218 382945 147454
rect 382597 147134 382945 147218
rect 382597 146898 382653 147134
rect 382889 146898 382945 147134
rect 382597 146866 382945 146898
rect 412863 147454 413211 147486
rect 412863 147218 412919 147454
rect 413155 147218 413211 147454
rect 412863 147134 413211 147218
rect 412863 146898 412919 147134
rect 413155 146898 413211 147134
rect 412863 146866 413211 146898
rect 506567 147454 506915 147486
rect 506567 147218 506623 147454
rect 506859 147218 506915 147454
rect 506567 147134 506915 147218
rect 506567 146898 506623 147134
rect 506859 146898 506915 147134
rect 506567 146866 506915 146898
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 289539 615218 289775 615454
rect 289539 614898 289775 615134
rect 505927 615218 506163 615454
rect 505927 614898 506163 615134
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 288779 597218 289015 597454
rect 288779 596898 289015 597134
rect 293967 597218 294203 597454
rect 293967 596898 294203 597134
rect 389031 597218 389267 597454
rect 389031 596898 389267 597134
rect 406395 597218 406631 597454
rect 406395 596898 406631 597134
rect 501459 597218 501695 597454
rect 501459 596898 501695 597134
rect 506687 597218 506923 597454
rect 506687 596898 506923 597134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 289539 579218 289775 579454
rect 289539 578898 289775 579134
rect 294647 579218 294883 579454
rect 294647 578898 294883 579134
rect 388351 579218 388587 579454
rect 388351 578898 388587 579134
rect 407075 579218 407311 579454
rect 407075 578898 407311 579134
rect 500779 579218 501015 579454
rect 500779 578898 501015 579134
rect 505927 579218 506163 579454
rect 505927 578898 506163 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 288779 561218 289015 561454
rect 288779 560898 289015 561134
rect 293967 561218 294203 561454
rect 293967 560898 294203 561134
rect 389031 561218 389267 561454
rect 389031 560898 389267 561134
rect 406395 561218 406631 561454
rect 406395 560898 406631 561134
rect 501459 561218 501695 561454
rect 501459 560898 501695 561134
rect 506687 561218 506923 561454
rect 506687 560898 506923 561134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 289539 543218 289775 543454
rect 289539 542898 289775 543134
rect 294647 543218 294883 543454
rect 294647 542898 294883 543134
rect 388351 543218 388587 543454
rect 388351 542898 388587 543134
rect 407075 543218 407311 543454
rect 407075 542898 407311 543134
rect 500779 543218 501015 543454
rect 500779 542898 501015 543134
rect 505927 543218 506163 543454
rect 505927 542898 506163 543134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 288269 489218 288505 489454
rect 288269 488898 288505 489134
rect 383333 489218 383569 489454
rect 383333 488898 383569 489134
rect 412239 489218 412475 489454
rect 412239 488898 412475 489134
rect 507303 489218 507539 489454
rect 507303 488898 507539 489134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 288949 471218 289185 471454
rect 288949 470898 289185 471134
rect 382653 471218 382889 471454
rect 382653 470898 382889 471134
rect 412919 471218 413155 471454
rect 412919 470898 413155 471134
rect 506623 471218 506859 471454
rect 506623 470898 506859 471134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 288269 453218 288505 453454
rect 288269 452898 288505 453134
rect 383333 453218 383569 453454
rect 383333 452898 383569 453134
rect 412239 453218 412475 453454
rect 412239 452898 412475 453134
rect 507303 453218 507539 453454
rect 507303 452898 507539 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 288949 435218 289185 435454
rect 288949 434898 289185 435134
rect 382653 435218 382889 435454
rect 382653 434898 382889 435134
rect 412919 435218 413155 435454
rect 412919 434898 413155 435134
rect 506623 435218 506859 435454
rect 506623 434898 506859 435134
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 288949 399218 289185 399454
rect 288949 398898 289185 399134
rect 382653 399218 382889 399454
rect 382653 398898 382889 399134
rect 412919 399218 413155 399454
rect 412919 398898 413155 399134
rect 506623 399218 506859 399454
rect 506623 398898 506859 399134
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 288269 381218 288505 381454
rect 288269 380898 288505 381134
rect 383333 381218 383569 381454
rect 383333 380898 383569 381134
rect 412239 381218 412475 381454
rect 412239 380898 412475 381134
rect 507303 381218 507539 381454
rect 507303 380898 507539 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 288949 363218 289185 363454
rect 288949 362898 289185 363134
rect 382653 363218 382889 363454
rect 382653 362898 382889 363134
rect 412919 363218 413155 363454
rect 412919 362898 413155 363134
rect 506623 363218 506859 363454
rect 506623 362898 506859 363134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 288269 345218 288505 345454
rect 288269 344898 288505 345134
rect 383333 345218 383569 345454
rect 383333 344898 383569 345134
rect 412239 345218 412475 345454
rect 412239 344898 412475 345134
rect 507303 345218 507539 345454
rect 507303 344898 507539 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 288949 291218 289185 291454
rect 288949 290898 289185 291134
rect 382653 291218 382889 291454
rect 382653 290898 382889 291134
rect 412919 291218 413155 291454
rect 412919 290898 413155 291134
rect 506623 291218 506859 291454
rect 506623 290898 506859 291134
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 288269 273218 288505 273454
rect 288269 272898 288505 273134
rect 383333 273218 383569 273454
rect 383333 272898 383569 273134
rect 412239 273218 412475 273454
rect 412239 272898 412475 273134
rect 507303 273218 507539 273454
rect 507303 272898 507539 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 288949 255218 289185 255454
rect 288949 254898 289185 255134
rect 382653 255218 382889 255454
rect 382653 254898 382889 255134
rect 412919 255218 413155 255454
rect 412919 254898 413155 255134
rect 506623 255218 506859 255454
rect 506623 254898 506859 255134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 288269 237218 288505 237454
rect 288269 236898 288505 237134
rect 383333 237218 383569 237454
rect 383333 236898 383569 237134
rect 412239 237218 412475 237454
rect 412239 236898 412475 237134
rect 507303 237218 507539 237454
rect 507303 236898 507539 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 288269 201218 288505 201454
rect 288269 200898 288505 201134
rect 383333 201218 383569 201454
rect 383333 200898 383569 201134
rect 412239 201218 412475 201454
rect 412239 200898 412475 201134
rect 507303 201218 507539 201454
rect 507303 200898 507539 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 288949 183218 289185 183454
rect 288949 182898 289185 183134
rect 382653 183218 382889 183454
rect 382653 182898 382889 183134
rect 412919 183218 413155 183454
rect 412919 182898 413155 183134
rect 506623 183218 506859 183454
rect 506623 182898 506859 183134
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 288269 165218 288505 165454
rect 288269 164898 288505 165134
rect 383333 165218 383569 165454
rect 383333 164898 383569 165134
rect 412239 165218 412475 165454
rect 412239 164898 412475 165134
rect 507303 165218 507539 165454
rect 507303 164898 507539 165134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 288949 147218 289185 147454
rect 288949 146898 289185 147134
rect 382653 147218 382889 147454
rect 382653 146898 382889 147134
rect 412919 147218 413155 147454
rect 412919 146898 413155 147134
rect 506623 147218 506859 147454
rect 506623 146898 506859 147134
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 289539 615454
rect 289775 615218 505927 615454
rect 506163 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 289539 615134
rect 289775 614898 505927 615134
rect 506163 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 288779 597454
rect 289015 597218 293967 597454
rect 294203 597218 389031 597454
rect 389267 597218 406395 597454
rect 406631 597218 501459 597454
rect 501695 597218 506687 597454
rect 506923 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 288779 597134
rect 289015 596898 293967 597134
rect 294203 596898 389031 597134
rect 389267 596898 406395 597134
rect 406631 596898 501459 597134
rect 501695 596898 506687 597134
rect 506923 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 289539 579454
rect 289775 579218 294647 579454
rect 294883 579218 388351 579454
rect 388587 579218 407075 579454
rect 407311 579218 500779 579454
rect 501015 579218 505927 579454
rect 506163 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 289539 579134
rect 289775 578898 294647 579134
rect 294883 578898 388351 579134
rect 388587 578898 407075 579134
rect 407311 578898 500779 579134
rect 501015 578898 505927 579134
rect 506163 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 288779 561454
rect 289015 561218 293967 561454
rect 294203 561218 389031 561454
rect 389267 561218 406395 561454
rect 406631 561218 501459 561454
rect 501695 561218 506687 561454
rect 506923 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 288779 561134
rect 289015 560898 293967 561134
rect 294203 560898 389031 561134
rect 389267 560898 406395 561134
rect 406631 560898 501459 561134
rect 501695 560898 506687 561134
rect 506923 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 289539 543454
rect 289775 543218 294647 543454
rect 294883 543218 388351 543454
rect 388587 543218 407075 543454
rect 407311 543218 500779 543454
rect 501015 543218 505927 543454
rect 506163 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 289539 543134
rect 289775 542898 294647 543134
rect 294883 542898 388351 543134
rect 388587 542898 407075 543134
rect 407311 542898 500779 543134
rect 501015 542898 505927 543134
rect 506163 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 288269 489454
rect 288505 489218 383333 489454
rect 383569 489218 412239 489454
rect 412475 489218 507303 489454
rect 507539 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 288269 489134
rect 288505 488898 383333 489134
rect 383569 488898 412239 489134
rect 412475 488898 507303 489134
rect 507539 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 288949 471454
rect 289185 471218 382653 471454
rect 382889 471218 412919 471454
rect 413155 471218 506623 471454
rect 506859 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 288949 471134
rect 289185 470898 382653 471134
rect 382889 470898 412919 471134
rect 413155 470898 506623 471134
rect 506859 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 288269 453454
rect 288505 453218 383333 453454
rect 383569 453218 412239 453454
rect 412475 453218 507303 453454
rect 507539 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 288269 453134
rect 288505 452898 383333 453134
rect 383569 452898 412239 453134
rect 412475 452898 507303 453134
rect 507539 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 288949 435454
rect 289185 435218 382653 435454
rect 382889 435218 412919 435454
rect 413155 435218 506623 435454
rect 506859 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 288949 435134
rect 289185 434898 382653 435134
rect 382889 434898 412919 435134
rect 413155 434898 506623 435134
rect 506859 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 288949 399454
rect 289185 399218 382653 399454
rect 382889 399218 412919 399454
rect 413155 399218 506623 399454
rect 506859 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 288949 399134
rect 289185 398898 382653 399134
rect 382889 398898 412919 399134
rect 413155 398898 506623 399134
rect 506859 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 288269 381454
rect 288505 381218 383333 381454
rect 383569 381218 412239 381454
rect 412475 381218 507303 381454
rect 507539 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 288269 381134
rect 288505 380898 383333 381134
rect 383569 380898 412239 381134
rect 412475 380898 507303 381134
rect 507539 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 288949 363454
rect 289185 363218 382653 363454
rect 382889 363218 412919 363454
rect 413155 363218 506623 363454
rect 506859 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 288949 363134
rect 289185 362898 382653 363134
rect 382889 362898 412919 363134
rect 413155 362898 506623 363134
rect 506859 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 288269 345454
rect 288505 345218 383333 345454
rect 383569 345218 412239 345454
rect 412475 345218 507303 345454
rect 507539 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 288269 345134
rect 288505 344898 383333 345134
rect 383569 344898 412239 345134
rect 412475 344898 507303 345134
rect 507539 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 288949 291454
rect 289185 291218 382653 291454
rect 382889 291218 412919 291454
rect 413155 291218 506623 291454
rect 506859 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 288949 291134
rect 289185 290898 382653 291134
rect 382889 290898 412919 291134
rect 413155 290898 506623 291134
rect 506859 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 288269 273454
rect 288505 273218 383333 273454
rect 383569 273218 412239 273454
rect 412475 273218 507303 273454
rect 507539 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 288269 273134
rect 288505 272898 383333 273134
rect 383569 272898 412239 273134
rect 412475 272898 507303 273134
rect 507539 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 288949 255454
rect 289185 255218 382653 255454
rect 382889 255218 412919 255454
rect 413155 255218 506623 255454
rect 506859 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 288949 255134
rect 289185 254898 382653 255134
rect 382889 254898 412919 255134
rect 413155 254898 506623 255134
rect 506859 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 288269 237454
rect 288505 237218 383333 237454
rect 383569 237218 412239 237454
rect 412475 237218 507303 237454
rect 507539 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 288269 237134
rect 288505 236898 383333 237134
rect 383569 236898 412239 237134
rect 412475 236898 507303 237134
rect 507539 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 288269 201454
rect 288505 201218 383333 201454
rect 383569 201218 412239 201454
rect 412475 201218 507303 201454
rect 507539 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 288269 201134
rect 288505 200898 383333 201134
rect 383569 200898 412239 201134
rect 412475 200898 507303 201134
rect 507539 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 288949 183454
rect 289185 183218 382653 183454
rect 382889 183218 412919 183454
rect 413155 183218 506623 183454
rect 506859 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 288949 183134
rect 289185 182898 382653 183134
rect 382889 182898 412919 183134
rect 413155 182898 506623 183134
rect 506859 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 288269 165454
rect 288505 165218 383333 165454
rect 383569 165218 412239 165454
rect 412475 165218 507303 165454
rect 507539 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 288269 165134
rect 288505 164898 383333 165134
rect 383569 164898 412239 165134
rect 412475 164898 507303 165134
rect 507539 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 288949 147454
rect 289185 147218 382653 147454
rect 382889 147218 412919 147454
rect 413155 147218 506623 147454
rect 506859 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 288949 147134
rect 289185 146898 382653 147134
rect 382889 146898 412919 147134
rect 413155 146898 506623 147134
rect 506859 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rest_top  mprj
timestamp 1640103014
transform 1 0 72000 0 1 60000
box 0 0 445188 579020
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 641020 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 641020 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 641020 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 641020 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 641020 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 641020 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 641020 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 641020 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 641020 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 641020 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 641020 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 641020 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 641020 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 641020 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 641020 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 641020 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 641020 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 641020 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 641020 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 641020 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 641020 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 641020 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 641020 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 641020 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 641020 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 641020 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 641020 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 641020 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 641020 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 641020 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 641020 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 641020 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 641020 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 641020 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 641020 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 641020 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 641020 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 641020 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 641020 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 641020 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 641020 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 641020 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 641020 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 641020 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 641020 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 641020 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 641020 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 641020 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 641020 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 641020 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 641020 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 641020 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 641020 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 641020 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 641020 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 641020 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 641020 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 641020 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 641020 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 641020 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 641020 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 641020 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 641020 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 641020 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 641020 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 641020 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 641020 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 641020 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 641020 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 641020 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 641020 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 641020 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 641020 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 641020 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 641020 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 641020 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 641020 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 641020 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 641020 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 641020 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 641020 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 641020 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 641020 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 641020 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 641020 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 641020 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 641020 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 641020 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 641020 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 641020 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 641020 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 641020 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 641020 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 641020 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 641020 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 641020 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 641020 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 641020 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 641020 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 641020 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
