magic
tech sky130A
timestamp 1640995782
<< nwell >>
rect -57 79 50 163
<< nmos >>
rect -11 2 4 44
<< pmos >>
rect -11 97 4 139
<< ndiff >>
rect -39 31 -11 44
rect -39 14 -34 31
rect -17 14 -11 31
rect -39 2 -11 14
rect 4 31 32 44
rect 4 14 10 31
rect 27 14 32 31
rect 4 2 32 14
<< pdiff >>
rect -39 127 -11 139
rect -39 110 -34 127
rect -17 110 -11 127
rect -39 97 -11 110
rect 4 127 32 139
rect 4 110 10 127
rect 27 110 32 127
rect 4 97 32 110
<< ndiffc >>
rect -34 14 -17 31
rect 10 14 27 31
<< pdiffc >>
rect -34 110 -17 127
rect 10 110 27 127
<< poly >>
rect -23 185 16 190
rect -23 168 -13 185
rect 6 168 16 185
rect -23 147 16 168
rect -11 139 4 147
rect -11 44 4 97
rect -11 -6 4 2
rect -23 -20 16 -6
rect -23 -37 -13 -20
rect 6 -37 16 -20
rect -23 -42 16 -37
<< polycont >>
rect -13 168 6 185
rect -13 -37 6 -20
<< locali >>
rect -23 185 16 190
rect -23 168 -13 185
rect 6 168 16 185
rect -23 156 16 168
rect -39 129 -13 139
rect -61 127 -13 129
rect -61 110 -34 127
rect -17 110 -13 127
rect -39 97 -13 110
rect 6 127 32 139
rect 6 110 10 127
rect 27 110 32 127
rect 6 97 32 110
rect 12 78 32 97
rect 12 58 43 78
rect 12 44 32 58
rect -39 31 -13 44
rect -59 14 -34 31
rect -17 14 -13 31
rect -59 12 -13 14
rect -39 2 -13 12
rect 6 31 32 44
rect 6 14 10 31
rect 27 14 32 31
rect 6 2 32 14
rect -23 -20 16 -15
rect -23 -37 -13 -20
rect 6 -37 16 -20
rect -23 -42 16 -37
<< viali >>
rect -13 168 6 185
rect -34 110 -17 127
rect -34 14 -17 31
rect -13 -37 6 -20
<< metal1 >>
rect -24 185 16 190
rect -24 168 -13 185
rect 6 168 16 185
rect -24 162 16 168
rect -40 127 -11 139
rect -40 110 -34 127
rect -17 110 -11 127
rect -40 97 -11 110
rect -39 31 -10 44
rect -39 14 -34 31
rect -17 14 -10 31
rect -39 2 -10 14
rect -24 -20 16 -14
rect -24 -37 -13 -20
rect 6 -37 16 -20
rect -24 -42 16 -37
<< end >>
