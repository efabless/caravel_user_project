magic
tech sky130A
magscale 1 2
timestamp 1640488860
<< poly >>
rect 1178 1088 1268 1098
rect 1178 1038 1198 1088
rect 1248 1038 1268 1088
rect 1178 1028 1268 1038
<< polycont >>
rect 1198 1038 1248 1088
<< locali >>
rect 1178 1088 1268 1098
rect 1178 1038 1198 1088
rect 1248 1038 1268 1088
rect 1178 1028 1268 1038
<< viali >>
rect 1198 1038 1248 1088
rect 3242 618 3282 664
rect 4876 624 4914 670
rect 1718 432 1758 478
rect 2030 470 2076 524
rect 3356 436 3394 488
rect 3662 476 3708 526
<< metal1 >>
rect 1536 1162 2002 1232
rect 1178 1088 1268 1098
rect 1178 1038 1198 1088
rect 1248 1048 1604 1088
rect 1248 1038 1268 1048
rect 1178 1028 1268 1038
rect 1552 780 1604 1048
rect 1916 914 2002 1162
rect 1552 742 3106 780
rect 1368 672 2094 712
rect 2026 558 2094 672
rect 2004 524 2096 558
rect 1696 478 1768 524
rect 1414 438 1718 478
rect 1414 312 1452 438
rect 1696 432 1718 438
rect 1758 432 1768 478
rect 2004 470 2030 524
rect 2076 470 2096 524
rect 3070 510 3106 742
rect 3232 688 3298 708
rect 4866 692 4924 714
rect 3232 664 3716 688
rect 3232 618 3242 664
rect 3282 652 3716 664
rect 3282 618 3298 652
rect 3232 576 3298 618
rect 3664 560 3716 652
rect 4866 670 4960 692
rect 4866 624 4876 670
rect 4914 654 4960 670
rect 4914 624 4924 654
rect 4866 570 4924 624
rect 3636 526 3742 560
rect 3342 510 3406 526
rect 3070 488 3406 510
rect 3070 474 3356 488
rect 2004 442 2096 470
rect 1696 368 1768 432
rect 3342 436 3356 474
rect 3394 436 3406 488
rect 3636 476 3662 526
rect 3708 476 3742 526
rect 3636 442 3742 476
rect 3342 390 3406 436
rect 452 272 1452 312
rect 1934 52 2020 166
rect 1598 -18 2020 52
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_1 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640415294
transform 1 0 3312 0 1 200
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_0
timestamp 1640415294
transform 1 0 1680 0 1 200
box -38 -49 1670 715
use doubletaillatchcomparator  doubletaillatchcomparator_0
timestamp 1640473169
transform 1 0 488 0 1 202
box -540 -220 1140 1030
<< labels >>
rlabel metal1 4960 674 4960 674 3 out
<< end >>
