magic
tech sky130A
timestamp 1640503333
<< nwell >>
rect -265 250 356 398
<< nmos >>
rect -200 40 -185 140
rect -135 40 -120 140
rect 0 40 15 140
rect 65 40 80 140
rect 150 40 165 140
rect 215 40 230 140
rect 280 40 295 140
rect 345 40 360 140
<< pmos >>
rect -200 275 -185 375
rect -135 275 -120 375
rect 0 275 15 375
rect 65 275 80 375
rect 150 275 165 375
rect 215 275 230 375
<< ndiff >>
rect -245 130 -200 140
rect -245 110 -235 130
rect -215 110 -200 130
rect -245 70 -200 110
rect -245 50 -235 70
rect -215 50 -200 70
rect -245 40 -200 50
rect -185 130 -135 140
rect -185 110 -170 130
rect -150 110 -135 130
rect -185 70 -135 110
rect -185 50 -170 70
rect -150 50 -135 70
rect -185 40 -135 50
rect -120 130 -75 140
rect -120 110 -105 130
rect -85 110 -75 130
rect -120 70 -75 110
rect -120 50 -105 70
rect -85 50 -75 70
rect -120 40 -75 50
rect -45 130 0 140
rect -45 110 -35 130
rect -15 110 0 130
rect -45 70 0 110
rect -45 50 -35 70
rect -15 50 0 70
rect -45 40 0 50
rect 15 130 65 140
rect 15 110 30 130
rect 50 110 65 130
rect 15 70 65 110
rect 15 50 30 70
rect 50 50 65 70
rect 15 40 65 50
rect 80 130 150 140
rect 80 110 105 130
rect 125 110 150 130
rect 80 70 150 110
rect 80 50 105 70
rect 125 50 150 70
rect 80 40 150 50
rect 165 130 215 140
rect 165 110 180 130
rect 200 110 215 130
rect 165 70 215 110
rect 165 50 180 70
rect 200 50 215 70
rect 165 40 215 50
rect 230 130 280 140
rect 230 110 245 130
rect 265 110 280 130
rect 230 70 280 110
rect 230 50 245 70
rect 265 50 280 70
rect 230 40 280 50
rect 295 130 345 140
rect 295 110 310 130
rect 330 110 345 130
rect 295 70 345 110
rect 295 50 310 70
rect 330 50 345 70
rect 295 40 345 50
rect 360 130 405 140
rect 360 110 375 130
rect 395 110 405 130
rect 360 70 405 110
rect 360 50 375 70
rect 395 50 405 70
rect 360 40 405 50
<< pdiff >>
rect -245 365 -200 375
rect -245 345 -235 365
rect -215 345 -200 365
rect -245 305 -200 345
rect -245 285 -235 305
rect -215 285 -200 305
rect -245 275 -200 285
rect -185 365 -135 375
rect -185 345 -170 365
rect -150 345 -135 365
rect -185 305 -135 345
rect -185 285 -170 305
rect -150 285 -135 305
rect -185 275 -135 285
rect -120 365 -75 375
rect -120 345 -105 365
rect -85 345 -75 365
rect -120 305 -75 345
rect -120 285 -105 305
rect -85 285 -75 305
rect -120 275 -75 285
rect -45 365 0 375
rect -45 345 -35 365
rect -15 345 0 365
rect -45 305 0 345
rect -45 285 -35 305
rect -15 285 0 305
rect -45 275 0 285
rect 15 365 65 375
rect 15 345 30 365
rect 50 345 65 365
rect 15 305 65 345
rect 15 285 30 305
rect 50 285 65 305
rect 15 275 65 285
rect 80 365 150 375
rect 80 345 105 365
rect 125 345 150 365
rect 80 305 150 345
rect 80 285 105 305
rect 125 285 150 305
rect 80 275 150 285
rect 165 365 215 375
rect 165 345 180 365
rect 200 345 215 365
rect 165 305 215 345
rect 165 285 180 305
rect 200 285 215 305
rect 165 275 215 285
rect 230 365 275 375
rect 230 345 245 365
rect 265 345 275 365
rect 230 305 275 345
rect 230 285 245 305
rect 265 285 275 305
rect 230 275 275 285
<< ndiffc >>
rect -235 110 -215 130
rect -235 50 -215 70
rect -170 110 -150 130
rect -170 50 -150 70
rect -105 110 -85 130
rect -105 50 -85 70
rect -35 110 -15 130
rect -35 50 -15 70
rect 30 110 50 130
rect 30 50 50 70
rect 105 110 125 130
rect 105 50 125 70
rect 180 110 200 130
rect 180 50 200 70
rect 245 110 265 130
rect 245 50 265 70
rect 310 110 330 130
rect 310 50 330 70
rect 375 110 395 130
rect 375 50 395 70
<< pdiffc >>
rect -235 345 -215 365
rect -235 285 -215 305
rect -170 345 -150 365
rect -170 285 -150 305
rect -105 345 -85 365
rect -105 285 -85 305
rect -35 345 -15 365
rect -35 285 -15 305
rect 30 345 50 365
rect 30 285 50 305
rect 105 345 125 365
rect 105 285 125 305
rect 180 345 200 365
rect 180 285 200 305
rect 245 345 265 365
rect 245 285 265 305
<< psubdiff >>
rect 460 -25 525 -15
rect 460 -60 475 -25
rect 510 -60 525 -25
rect 460 -70 525 -60
<< nsubdiff >>
rect 275 360 335 375
rect 275 340 305 360
rect 325 340 335 360
rect 275 320 335 340
rect 275 300 305 320
rect 325 300 335 320
rect 275 275 335 300
<< psubdiffcont >>
rect 475 -60 510 -25
<< nsubdiffcont >>
rect 305 340 325 360
rect 305 300 325 320
<< poly >>
rect -200 465 360 480
rect -200 430 -185 465
rect -230 425 -185 430
rect -230 400 -220 425
rect -195 405 -185 425
rect -70 435 -25 440
rect -70 410 -60 435
rect -35 430 -25 435
rect -35 415 230 430
rect -35 410 -25 415
rect -70 405 -25 410
rect -195 400 -120 405
rect -230 395 -120 400
rect -200 390 -120 395
rect -200 375 -185 390
rect -135 375 -120 390
rect 0 375 15 390
rect 65 375 80 390
rect 150 375 165 390
rect 215 375 230 415
rect -200 260 -185 275
rect -135 260 -120 275
rect 0 235 15 275
rect -245 230 15 235
rect -245 205 -235 230
rect -210 220 15 230
rect 65 255 80 275
rect 65 250 110 255
rect 65 225 75 250
rect 100 225 110 250
rect 65 220 110 225
rect -210 205 -200 220
rect -245 200 -200 205
rect -200 140 -185 155
rect -135 140 -120 155
rect 0 140 15 155
rect 65 140 80 220
rect 150 195 165 275
rect 215 260 230 275
rect 120 190 165 195
rect 120 165 130 190
rect 155 165 165 190
rect 120 160 165 165
rect 150 140 165 160
rect 215 140 230 155
rect 280 140 295 155
rect 345 140 360 465
rect -200 15 -185 40
rect -230 10 -185 15
rect -230 -15 -220 10
rect -195 -15 -185 10
rect -135 15 -120 40
rect -135 10 -75 15
rect -135 0 -110 10
rect -230 -20 -185 -15
rect -120 -15 -110 0
rect -85 -15 -75 10
rect -120 -20 -75 -15
rect 0 0 15 40
rect 65 25 80 40
rect 150 25 165 40
rect 215 0 230 40
rect 280 0 295 40
rect 345 25 360 40
rect 0 -15 295 0
rect 0 -20 35 -15
rect -10 -30 35 -20
rect -10 -55 0 -30
rect 25 -55 35 -30
rect -10 -60 35 -55
<< polycont >>
rect -220 400 -195 425
rect -60 410 -35 435
rect -235 205 -210 230
rect 75 225 100 250
rect 130 165 155 190
rect -220 -15 -195 10
rect -110 -15 -85 10
rect 0 -55 25 -30
<< locali >>
rect -180 490 -130 500
rect -180 460 -170 490
rect -140 460 -130 490
rect -180 450 -130 460
rect 90 490 140 500
rect 90 460 100 490
rect 130 460 140 490
rect 90 450 140 460
rect -230 425 -185 430
rect -230 400 -220 425
rect -195 400 -185 425
rect -230 395 -185 400
rect -165 375 -145 450
rect -70 435 -25 440
rect -70 425 -60 435
rect -95 410 -60 425
rect -35 410 -25 435
rect -95 405 -25 410
rect 105 415 125 450
rect -95 375 -75 405
rect 105 395 315 415
rect 105 375 125 395
rect -245 365 -205 375
rect -245 345 -235 365
rect -215 345 -205 365
rect -245 305 -205 345
rect -245 285 -235 305
rect -215 285 -205 305
rect -245 275 -205 285
rect -180 365 -140 375
rect -180 345 -170 365
rect -150 345 -140 365
rect -180 305 -140 345
rect -180 285 -170 305
rect -150 285 -140 305
rect -180 275 -140 285
rect -115 365 -75 375
rect -115 345 -105 365
rect -85 345 -75 365
rect -115 305 -75 345
rect -115 285 -105 305
rect -85 285 -75 305
rect -115 275 -75 285
rect -45 365 -5 375
rect -45 345 -35 365
rect -15 345 -5 365
rect -45 305 -5 345
rect -45 285 -35 305
rect -15 285 -5 305
rect -45 275 -5 285
rect 20 365 60 375
rect 20 345 30 365
rect 50 345 60 365
rect 20 305 60 345
rect 20 285 30 305
rect 50 285 60 305
rect 20 275 60 285
rect 95 365 135 375
rect 95 345 105 365
rect 125 345 135 365
rect 95 305 135 345
rect 95 285 105 305
rect 125 285 135 305
rect 95 275 135 285
rect 170 365 210 375
rect 170 345 180 365
rect 200 345 210 365
rect 170 305 210 345
rect 170 285 180 305
rect 200 285 210 305
rect 170 275 210 285
rect 235 365 275 375
rect 235 345 245 365
rect 265 345 275 365
rect 235 305 275 345
rect 235 285 245 305
rect 265 285 275 305
rect 295 365 315 395
rect 295 360 335 365
rect 295 340 305 360
rect 325 340 335 360
rect 295 320 335 340
rect 295 300 305 320
rect 325 300 335 320
rect 295 290 335 300
rect 235 275 275 285
rect -245 235 -225 275
rect -245 230 -200 235
rect -245 205 -235 230
rect -210 205 -200 230
rect -245 200 -200 205
rect -245 140 -225 200
rect -95 140 -75 275
rect -35 180 -15 275
rect 250 255 270 275
rect 65 250 270 255
rect 65 225 75 250
rect 100 235 270 250
rect 100 225 110 235
rect 65 220 110 225
rect 120 190 165 195
rect 120 180 130 190
rect -35 165 130 180
rect 155 165 165 190
rect -35 160 165 165
rect 25 140 45 160
rect 185 140 205 235
rect 320 160 525 180
rect 320 140 340 160
rect -245 130 -205 140
rect -245 110 -235 130
rect -215 110 -205 130
rect -245 70 -205 110
rect -245 50 -235 70
rect -215 50 -205 70
rect -245 40 -205 50
rect -180 130 -140 140
rect -180 110 -170 130
rect -150 110 -140 130
rect -180 70 -140 110
rect -180 50 -170 70
rect -150 50 -140 70
rect -180 40 -140 50
rect -115 130 -75 140
rect -115 110 -105 130
rect -85 110 -75 130
rect -115 70 -75 110
rect -115 50 -105 70
rect -85 50 -75 70
rect -115 40 -75 50
rect -45 130 -5 140
rect -45 110 -35 130
rect -15 110 -5 130
rect -45 70 -5 110
rect -45 50 -35 70
rect -15 50 -5 70
rect -45 40 -5 50
rect 20 130 60 140
rect 20 110 30 130
rect 50 110 60 130
rect 20 70 60 110
rect 20 50 30 70
rect 50 50 60 70
rect 20 40 60 50
rect 95 130 135 140
rect 95 110 105 130
rect 125 110 135 130
rect 95 70 135 110
rect 95 50 105 70
rect 125 50 135 70
rect 95 40 135 50
rect 170 130 210 140
rect 170 110 180 130
rect 200 110 210 130
rect 170 70 210 110
rect 170 50 180 70
rect 200 50 210 70
rect 170 40 210 50
rect 235 130 275 140
rect 235 110 245 130
rect 265 110 275 130
rect 235 70 275 110
rect 235 50 245 70
rect 265 50 275 70
rect 235 40 275 50
rect 300 130 340 140
rect 300 110 310 130
rect 330 110 340 130
rect 300 70 340 110
rect 300 50 310 70
rect 330 50 340 70
rect 300 40 340 50
rect 365 130 405 140
rect 365 110 375 130
rect 395 110 405 130
rect 365 70 405 110
rect 365 50 375 70
rect 395 50 405 70
rect 365 40 405 50
rect 505 100 525 160
rect 505 90 560 100
rect 505 55 515 90
rect 550 55 560 90
rect 505 45 560 55
rect -230 10 -185 15
rect -230 -15 -220 10
rect -195 -15 -185 10
rect -230 -20 -185 -15
rect -165 -80 -145 40
rect -45 20 -25 40
rect 105 20 125 40
rect 255 20 275 40
rect -45 15 275 20
rect -120 10 -75 15
rect -120 -15 -110 10
rect -85 -15 -75 10
rect -45 0 175 15
rect 165 -5 175 0
rect 195 0 275 15
rect 195 -5 205 0
rect 165 -10 205 -5
rect -120 -20 -75 -15
rect 385 -20 405 40
rect -10 -30 35 -20
rect -10 -55 0 -30
rect 25 -55 35 -30
rect -10 -60 35 -55
rect 360 -40 405 -20
rect 460 -25 525 -15
rect 360 -80 380 -40
rect 460 -60 475 -25
rect 510 -60 525 -25
rect -165 -100 380 -80
rect 460 -70 525 -60
<< viali >>
rect -170 460 -140 490
rect 100 460 130 490
rect -220 400 -195 425
rect 130 165 155 190
rect 515 55 550 90
rect -220 -15 -195 10
rect -110 -15 -85 10
rect 175 -5 195 15
rect 0 -55 25 -30
rect 475 -60 510 -25
rect 405 -90 435 -60
<< metal1 >>
rect -270 490 570 515
rect -270 480 -170 490
rect -180 460 -170 480
rect -140 480 100 490
rect -140 460 -130 480
rect -180 450 -130 460
rect 90 460 100 480
rect 130 480 570 490
rect 130 460 140 480
rect 90 450 140 460
rect -270 425 -185 430
rect -270 410 -220 425
rect -230 400 -220 410
rect -195 400 -185 425
rect -230 395 -185 400
rect 120 190 570 195
rect 120 165 130 190
rect 155 175 570 190
rect 155 165 165 175
rect 120 160 165 165
rect 505 90 560 100
rect 505 55 515 90
rect 550 55 560 90
rect -270 35 10 55
rect 505 45 560 55
rect -230 10 -185 15
rect -230 0 -220 10
rect -270 -15 -220 0
rect -195 -15 -185 10
rect -270 -20 -185 -15
rect -120 10 -75 15
rect -120 -15 -110 10
rect -85 -15 -75 10
rect -120 -20 -75 -15
rect -10 -20 10 35
rect 165 15 205 20
rect 165 -5 175 15
rect 195 -5 205 15
rect 165 -10 205 -5
rect -120 -35 -100 -20
rect -270 -55 -100 -35
rect -10 -30 35 -20
rect -10 -55 0 -30
rect 25 -55 35 -30
rect -10 -60 35 -55
rect 175 -75 195 -10
rect 460 -25 525 -15
rect 460 -50 475 -25
rect 395 -60 475 -50
rect 510 -60 525 -25
rect 395 -75 405 -60
rect -270 -90 405 -75
rect 435 -75 525 -60
rect 435 -90 570 -75
rect -270 -110 570 -90
<< via1 >>
rect 515 55 550 90
rect 405 -90 435 -60
<< metal2 >>
rect 505 90 560 100
rect 505 55 515 90
rect 550 55 560 90
rect 505 45 560 55
rect 395 -60 445 -50
rect 395 -90 405 -60
rect 435 -90 445 -60
rect 395 -100 445 -90
<< via2 >>
rect 515 55 550 90
rect 405 -90 435 -60
<< metal3 >>
rect -240 -10 465 515
rect 505 90 560 100
rect 505 55 515 90
rect 550 55 560 90
rect 505 45 560 55
rect 415 -50 445 -10
rect 395 -60 445 -50
rect 395 -90 405 -60
rect 435 -90 445 -60
rect 395 -100 445 -90
<< via3 >>
rect 515 55 550 90
<< mimcap >>
rect -225 85 450 500
rect -225 50 405 85
rect 440 50 450 85
rect -225 5 450 50
<< mimcapcontact >>
rect 405 50 440 85
<< metal4 >>
rect 505 95 560 100
rect 400 90 560 95
rect 400 85 515 90
rect 400 50 405 85
rect 440 55 515 85
rect 550 55 560 90
rect 440 50 560 55
rect 400 45 560 50
<< labels >>
rlabel metal1 -270 -15 -270 -15 7 Vref1
rlabel metal1 -270 425 -270 425 7 clk
rlabel metal1 -270 -90 -270 -90 7 GND
rlabel metal1 -270 490 -270 490 7 VDD
rlabel metal1 -270 45 -270 45 7 clkbar
rlabel metal1 -270 -45 -270 -45 7 vref2
rlabel metal1 569 -95 570 -95 3 gnd
rlabel metal1 569 497 570 497 3 vdd
rlabel metal1 570 186 570 186 3 out
<< end >>
