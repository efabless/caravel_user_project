VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_32x256_8
   CLASS BLOCK ;
   SIZE 475.7 BY 394.78 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.72 0.0 105.1 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 0.0 111.22 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.08 0.0 123.46 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.52 0.0 128.9 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.96 0.0 134.34 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 0.0 146.58 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 0.0 152.02 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 0.0 157.46 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  175.44 0.0 175.82 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 0.0 181.26 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 0.0 186.7 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 0.0 199.62 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 0.0 205.06 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.62 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  251.6 0.0 251.98 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 0.0 268.3 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 0.0 281.22 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 0.0 286.66 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.48 0.0 75.86 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 127.16 0.38 127.54 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 135.32 0.38 135.7 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.76 0.38 141.14 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.92 0.38 149.3 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.36 0.38 154.74 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.2 0.38 163.58 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 0.38 169.02 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  395.08 394.4 395.46 394.78 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  475.32 81.6 475.7 81.98 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  475.32 73.44 475.7 73.82 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  475.32 67.32 475.7 67.7 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  413.44 0.0 413.82 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  411.4 0.0 411.78 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  412.08 0.0 412.46 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  412.76 0.0 413.14 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 25.16 0.38 25.54 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  475.32 381.48 475.7 381.86 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 34.0 0.38 34.38 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  27.2 0.0 27.58 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  448.12 394.4 448.5 394.78 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  81.6 0.0 81.98 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.04 0.0 87.42 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 0.0 94.22 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.6 0.0 98.98 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.36 0.0 137.74 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 0.0 144.54 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.6 0.0 149.98 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 0.0 164.26 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 0.0 170.38 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 0.0 182.62 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.0 0.0 187.38 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 0.0 194.86 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 0.0 207.78 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.52 0.0 213.9 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.76 0.0 226.14 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.2 0.0 231.58 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  237.32 0.0 237.7 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.84 0.0 264.22 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 0.0 270.34 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 0.0 282.58 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.96 0.0 287.34 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 0.0 294.82 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 0.0 300.94 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 0.0 307.74 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  313.48 0.0 313.86 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 0.0 319.98 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 0.0 326.1 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.84 0.0 332.22 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  138.72 394.4 139.1 394.78 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  145.52 394.4 145.9 394.78 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 394.4 151.34 394.78 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 394.4 158.14 394.78 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 394.4 164.26 394.78 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 394.4 171.06 394.78 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 394.4 177.18 394.78 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 394.4 182.62 394.78 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 394.4 189.42 394.78 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 394.4 194.86 394.78 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 394.4 201.66 394.78 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 394.4 207.78 394.78 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 394.4 214.58 394.78 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 394.4 220.02 394.78 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.76 394.4 226.14 394.78 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 394.4 232.94 394.78 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 394.4 239.06 394.78 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 394.4 245.86 394.78 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 394.4 251.3 394.78 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 394.4 258.1 394.78 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 394.4 263.54 394.78 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 394.4 269.66 394.78 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 394.4 276.46 394.78 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 394.4 282.58 394.78 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 394.4 289.38 394.78 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 394.4 294.82 394.78 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 394.4 301.62 394.78 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 394.4 307.74 394.78 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  314.16 394.4 314.54 394.78 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  319.6 394.4 319.98 394.78 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 394.4 326.1 394.78 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  332.52 394.4 332.9 394.78 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  1.36 391.68 474.34 393.42 ;
         LAYER met4 ;
         RECT  472.6 1.36 474.34 393.42 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 393.42 ;
         LAYER met3 ;
         RECT  1.36 1.36 474.34 3.1 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 388.28 470.94 390.02 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 390.02 ;
         LAYER met3 ;
         RECT  4.76 4.76 470.94 6.5 ;
         LAYER met4 ;
         RECT  469.2 4.76 470.94 390.02 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 475.08 394.16 ;
   LAYER  met2 ;
      RECT  0.62 0.62 475.08 394.16 ;
   LAYER  met3 ;
      RECT  0.98 126.56 475.08 128.14 ;
      RECT  0.62 128.14 0.98 134.72 ;
      RECT  0.62 136.3 0.98 140.16 ;
      RECT  0.62 141.74 0.98 148.32 ;
      RECT  0.62 149.9 0.98 153.76 ;
      RECT  0.62 155.34 0.98 162.6 ;
      RECT  0.62 164.18 0.98 168.04 ;
      RECT  0.98 81.0 474.72 82.58 ;
      RECT  0.98 82.58 474.72 126.56 ;
      RECT  474.72 82.58 475.08 126.56 ;
      RECT  474.72 74.42 475.08 81.0 ;
      RECT  474.72 68.3 475.08 72.84 ;
      RECT  0.98 128.14 474.72 380.88 ;
      RECT  0.98 380.88 474.72 382.46 ;
      RECT  474.72 128.14 475.08 380.88 ;
      RECT  0.62 26.14 0.98 33.4 ;
      RECT  0.62 34.98 0.98 126.56 ;
      RECT  0.62 169.62 0.76 391.08 ;
      RECT  0.62 391.08 0.76 394.02 ;
      RECT  0.62 394.02 0.76 394.16 ;
      RECT  0.76 169.62 0.98 391.08 ;
      RECT  0.76 394.02 0.98 394.16 ;
      RECT  0.98 394.02 474.72 394.16 ;
      RECT  474.72 382.46 474.94 391.08 ;
      RECT  474.72 394.02 474.94 394.16 ;
      RECT  474.94 382.46 475.08 391.08 ;
      RECT  474.94 391.08 475.08 394.02 ;
      RECT  474.94 394.02 475.08 394.16 ;
      RECT  0.98 0.62 474.72 0.76 ;
      RECT  474.72 0.62 474.94 0.76 ;
      RECT  474.72 3.7 474.94 66.72 ;
      RECT  474.94 0.62 475.08 0.76 ;
      RECT  474.94 0.76 475.08 3.7 ;
      RECT  474.94 3.7 475.08 66.72 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 24.56 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 24.56 ;
      RECT  0.98 382.46 4.16 387.68 ;
      RECT  0.98 387.68 4.16 390.62 ;
      RECT  0.98 390.62 4.16 391.08 ;
      RECT  4.16 382.46 471.54 387.68 ;
      RECT  4.16 390.62 471.54 391.08 ;
      RECT  471.54 382.46 474.72 387.68 ;
      RECT  471.54 387.68 474.72 390.62 ;
      RECT  471.54 390.62 474.72 391.08 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 81.0 ;
      RECT  4.16 3.7 471.54 4.16 ;
      RECT  4.16 7.1 471.54 81.0 ;
      RECT  471.54 3.7 474.72 4.16 ;
      RECT  471.54 4.16 474.72 7.1 ;
      RECT  471.54 7.1 474.72 81.0 ;
   LAYER  met4 ;
      RECT  104.12 0.98 105.7 394.16 ;
      RECT  105.7 0.62 110.24 0.98 ;
      RECT  111.82 0.62 115.68 0.98 ;
      RECT  117.26 0.62 122.48 0.98 ;
      RECT  124.06 0.62 127.92 0.98 ;
      RECT  129.5 0.62 133.36 0.98 ;
      RECT  152.62 0.62 156.48 0.98 ;
      RECT  258.02 0.62 261.88 0.98 ;
      RECT  105.7 0.98 394.48 393.8 ;
      RECT  394.48 0.98 396.06 393.8 ;
      RECT  28.18 0.62 74.88 0.98 ;
      RECT  396.06 393.8 447.52 394.16 ;
      RECT  76.46 0.62 81.0 0.98 ;
      RECT  82.58 0.62 86.44 0.98 ;
      RECT  88.02 0.62 93.24 0.98 ;
      RECT  94.82 0.62 98.0 0.98 ;
      RECT  99.58 0.62 104.12 0.98 ;
      RECT  134.94 0.62 136.76 0.98 ;
      RECT  138.34 0.62 138.8 0.98 ;
      RECT  140.38 0.62 143.56 0.98 ;
      RECT  145.14 0.62 145.6 0.98 ;
      RECT  147.18 0.62 149.0 0.98 ;
      RECT  150.58 0.62 151.04 0.98 ;
      RECT  158.74 0.62 162.6 0.98 ;
      RECT  164.86 0.62 168.04 0.98 ;
      RECT  170.98 0.62 174.84 0.98 ;
      RECT  177.1 0.62 180.28 0.98 ;
      RECT  183.22 0.62 185.72 0.98 ;
      RECT  187.98 0.62 191.84 0.98 ;
      RECT  193.42 0.62 193.88 0.98 ;
      RECT  195.46 0.62 198.64 0.98 ;
      RECT  200.22 0.62 200.68 0.98 ;
      RECT  202.26 0.62 204.08 0.98 ;
      RECT  205.66 0.62 206.8 0.98 ;
      RECT  208.38 0.62 209.52 0.98 ;
      RECT  211.1 0.62 212.92 0.98 ;
      RECT  214.5 0.62 214.96 0.98 ;
      RECT  216.54 0.62 219.04 0.98 ;
      RECT  220.62 0.62 221.76 0.98 ;
      RECT  223.34 0.62 225.16 0.98 ;
      RECT  226.74 0.62 227.2 0.98 ;
      RECT  228.78 0.62 230.6 0.98 ;
      RECT  232.18 0.62 232.64 0.98 ;
      RECT  234.22 0.62 236.72 0.98 ;
      RECT  238.3 0.62 238.76 0.98 ;
      RECT  240.34 0.62 242.84 0.98 ;
      RECT  245.78 0.62 250.32 0.98 ;
      RECT  252.58 0.62 254.4 0.98 ;
      RECT  255.98 0.62 256.44 0.98 ;
      RECT  264.82 0.62 267.32 0.98 ;
      RECT  268.9 0.62 269.36 0.98 ;
      RECT  270.94 0.62 273.44 0.98 ;
      RECT  275.02 0.62 275.48 0.98 ;
      RECT  277.06 0.62 280.24 0.98 ;
      RECT  283.18 0.62 285.68 0.98 ;
      RECT  287.94 0.62 293.84 0.98 ;
      RECT  295.42 0.62 299.96 0.98 ;
      RECT  301.54 0.62 306.76 0.98 ;
      RECT  308.34 0.62 312.88 0.98 ;
      RECT  314.46 0.62 319.0 0.98 ;
      RECT  320.58 0.62 325.12 0.98 ;
      RECT  326.7 0.62 331.24 0.98 ;
      RECT  332.82 0.62 410.8 0.98 ;
      RECT  105.7 393.8 138.12 394.16 ;
      RECT  139.7 393.8 144.92 394.16 ;
      RECT  146.5 393.8 150.36 394.16 ;
      RECT  151.94 393.8 157.16 394.16 ;
      RECT  158.74 393.8 163.28 394.16 ;
      RECT  164.86 393.8 170.08 394.16 ;
      RECT  171.66 393.8 176.2 394.16 ;
      RECT  177.78 393.8 181.64 394.16 ;
      RECT  183.22 393.8 188.44 394.16 ;
      RECT  190.02 393.8 193.88 394.16 ;
      RECT  195.46 393.8 200.68 394.16 ;
      RECT  202.26 393.8 206.8 394.16 ;
      RECT  208.38 393.8 213.6 394.16 ;
      RECT  215.18 393.8 219.04 394.16 ;
      RECT  220.62 393.8 225.16 394.16 ;
      RECT  226.74 393.8 231.96 394.16 ;
      RECT  233.54 393.8 238.08 394.16 ;
      RECT  239.66 393.8 244.88 394.16 ;
      RECT  246.46 393.8 250.32 394.16 ;
      RECT  251.9 393.8 257.12 394.16 ;
      RECT  258.7 393.8 262.56 394.16 ;
      RECT  264.14 393.8 268.68 394.16 ;
      RECT  270.26 393.8 275.48 394.16 ;
      RECT  277.06 393.8 281.6 394.16 ;
      RECT  283.18 393.8 288.4 394.16 ;
      RECT  289.98 393.8 293.84 394.16 ;
      RECT  295.42 393.8 300.64 394.16 ;
      RECT  302.22 393.8 306.76 394.16 ;
      RECT  308.34 393.8 313.56 394.16 ;
      RECT  315.14 393.8 319.0 394.16 ;
      RECT  320.58 393.8 325.12 394.16 ;
      RECT  326.7 393.8 331.92 394.16 ;
      RECT  333.5 393.8 394.48 394.16 ;
      RECT  474.94 0.98 475.08 393.8 ;
      RECT  414.42 0.62 472.0 0.76 ;
      RECT  414.42 0.76 472.0 0.98 ;
      RECT  472.0 0.62 474.94 0.76 ;
      RECT  474.94 0.62 475.08 0.76 ;
      RECT  474.94 0.76 475.08 0.98 ;
      RECT  449.1 393.8 472.0 394.02 ;
      RECT  449.1 394.02 472.0 394.16 ;
      RECT  472.0 394.02 474.94 394.16 ;
      RECT  474.94 393.8 475.08 394.02 ;
      RECT  474.94 394.02 475.08 394.16 ;
      RECT  0.62 0.98 0.76 394.02 ;
      RECT  0.62 394.02 0.76 394.16 ;
      RECT  0.76 394.02 3.7 394.16 ;
      RECT  3.7 394.02 104.12 394.16 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 26.6 0.76 ;
      RECT  3.7 0.76 26.6 0.98 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 390.62 ;
      RECT  3.7 390.62 4.16 394.02 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 390.62 7.1 394.02 ;
      RECT  7.1 0.98 104.12 4.16 ;
      RECT  7.1 4.16 104.12 390.62 ;
      RECT  7.1 390.62 104.12 394.02 ;
      RECT  396.06 0.98 468.6 4.16 ;
      RECT  396.06 4.16 468.6 390.62 ;
      RECT  396.06 390.62 468.6 393.8 ;
      RECT  468.6 0.98 471.54 4.16 ;
      RECT  468.6 390.62 471.54 393.8 ;
      RECT  471.54 0.98 472.0 4.16 ;
      RECT  471.54 4.16 472.0 390.62 ;
      RECT  471.54 390.62 472.0 393.8 ;
   END
END    sky130_sram_1kbyte_1rw1r_32x256_8
END    LIBRARY
