magic
tech sky130A
timestamp 1641069145
<< nwell >>
rect -66 75 146 184
<< nmos >>
rect -3 -1 12 41
<< pmos >>
rect -3 94 12 136
<< ndiff >>
rect -31 28 -3 41
rect -31 11 -26 28
rect -9 11 -3 28
rect -31 -1 -3 11
rect 12 28 40 41
rect 12 11 18 28
rect 35 11 40 28
rect 12 -1 40 11
<< pdiff >>
rect -31 123 -3 136
rect -31 106 -26 123
rect -9 106 -3 123
rect -31 94 -3 106
rect 12 123 40 136
rect 12 106 18 123
rect 35 106 40 123
rect 12 94 40 106
<< ndiffc >>
rect -26 11 -9 28
rect 18 11 35 28
<< pdiffc >>
rect -26 106 -9 123
rect 18 106 35 123
<< poly >>
rect -15 177 24 184
rect -15 160 -5 177
rect 14 160 24 177
rect -15 144 24 160
rect -3 136 12 144
rect -3 41 12 94
rect -3 -9 12 -1
rect -15 -23 24 -9
rect -15 -40 -5 -23
rect 14 -40 24 -23
rect -15 -45 24 -40
<< polycont >>
rect -5 160 14 177
rect -5 -40 14 -23
<< locali >>
rect -54 177 -32 180
rect -54 160 -52 177
rect -35 160 -32 177
rect -54 158 -32 160
rect -50 136 -32 158
rect -15 177 24 184
rect -15 160 -5 177
rect 14 160 24 177
rect -15 153 24 160
rect -50 123 -5 136
rect -50 106 -26 123
rect -9 106 -5 123
rect -50 94 -5 106
rect 14 123 40 136
rect 14 106 18 123
rect 35 106 40 123
rect 14 94 40 106
rect 17 78 40 94
rect 17 61 20 78
rect 37 61 40 78
rect 17 58 40 61
rect -31 28 -5 41
rect -31 11 -26 28
rect -9 11 -5 28
rect -31 -1 -5 11
rect 14 28 40 41
rect 14 11 18 28
rect 35 11 40 28
rect 14 -1 40 11
rect -15 -23 24 -18
rect -15 -40 -5 -23
rect 14 -40 24 -23
rect -15 -45 24 -40
rect 59 -45 86 184
<< viali >>
rect -52 160 -35 177
rect 20 61 37 78
rect -26 11 -9 28
rect 18 11 35 28
<< metal1 >>
rect -66 179 -32 184
rect -66 177 146 179
rect -66 160 -52 177
rect -35 160 146 177
rect -66 159 146 160
rect -66 153 -32 159
rect 14 78 43 84
rect 14 77 20 78
rect -66 61 20 77
rect 37 77 43 78
rect 37 61 146 77
rect -66 57 146 61
rect -31 31 -3 34
rect 14 31 40 34
rect -66 28 -3 31
rect -66 11 -26 28
rect -9 11 -3 28
rect -66 9 -3 11
rect 12 28 146 31
rect 12 11 18 28
rect 35 11 146 28
rect 12 9 146 11
rect -31 5 -3 9
rect 14 5 40 9
<< end >>
