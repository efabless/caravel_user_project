magic
tech sky130A
magscale 1 2
timestamp 1640415294
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 214 229 959 273
rect 1443 229 1631 241
rect 214 180 1631 229
rect 1 49 1631 180
rect 0 0 1632 49
<< scnmos >>
rect 293 163 323 247
rect 424 163 454 247
rect 510 163 540 247
rect 596 163 626 247
rect 668 163 698 247
rect 80 70 110 154
rect 850 119 880 247
rect 948 119 978 203
rect 1086 119 1116 203
rect 1158 119 1188 203
rect 1259 75 1289 203
rect 1522 47 1552 215
<< scpmoshvt >>
rect 80 468 110 596
rect 270 413 300 541
rect 410 413 440 497
rect 496 413 526 497
rect 636 413 666 497
rect 708 413 738 497
rect 825 379 855 547
rect 927 379 957 547
rect 1086 379 1116 463
rect 1158 379 1188 463
rect 1267 379 1297 547
rect 1522 367 1552 619
<< ndiff >>
rect 240 221 293 247
rect 240 187 248 221
rect 282 187 293 221
rect 240 163 293 187
rect 323 205 424 247
rect 323 171 358 205
rect 392 171 424 205
rect 323 163 424 171
rect 454 222 510 247
rect 454 188 465 222
rect 499 188 510 222
rect 454 163 510 188
rect 540 222 596 247
rect 540 188 551 222
rect 585 188 596 222
rect 540 163 596 188
rect 626 163 668 247
rect 698 182 850 247
rect 698 163 730 182
rect 27 129 80 154
rect 27 95 35 129
rect 69 95 80 129
rect 27 70 80 95
rect 110 130 163 154
rect 110 96 121 130
rect 155 96 163 130
rect 110 70 163 96
rect 722 148 730 163
rect 764 148 798 182
rect 832 148 850 182
rect 722 119 850 148
rect 880 233 933 247
rect 880 199 891 233
rect 925 203 933 233
rect 1469 203 1522 215
rect 925 199 948 203
rect 880 165 948 199
rect 880 131 897 165
rect 931 131 948 165
rect 880 119 948 131
rect 978 178 1086 203
rect 978 144 1014 178
rect 1048 144 1086 178
rect 978 119 1086 144
rect 1116 119 1158 203
rect 1188 189 1259 203
rect 1188 155 1211 189
rect 1245 155 1259 189
rect 1188 121 1259 155
rect 1188 119 1211 121
rect 1203 87 1211 119
rect 1245 87 1259 121
rect 1203 75 1259 87
rect 1289 189 1353 203
rect 1289 155 1311 189
rect 1345 155 1353 189
rect 1289 121 1353 155
rect 1289 87 1311 121
rect 1345 87 1353 121
rect 1289 75 1353 87
rect 1469 169 1477 203
rect 1511 169 1522 203
rect 1469 93 1522 169
rect 1469 59 1477 93
rect 1511 59 1522 93
rect 1469 47 1522 59
rect 1552 203 1605 215
rect 1552 169 1563 203
rect 1597 169 1605 203
rect 1552 101 1605 169
rect 1552 67 1563 101
rect 1597 67 1605 101
rect 1552 47 1605 67
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 515 80 550
rect 27 481 35 515
rect 69 481 80 515
rect 27 468 80 481
rect 110 582 163 596
rect 110 548 121 582
rect 155 548 163 582
rect 110 514 163 548
rect 110 480 121 514
rect 155 480 163 514
rect 110 468 163 480
rect 217 527 270 541
rect 217 493 225 527
rect 259 493 270 527
rect 217 459 270 493
rect 217 425 225 459
rect 259 425 270 459
rect 217 413 270 425
rect 300 510 353 541
rect 300 476 311 510
rect 345 497 353 510
rect 760 561 810 573
rect 760 527 768 561
rect 802 547 810 561
rect 1469 607 1522 619
rect 1469 573 1477 607
rect 1511 573 1522 607
rect 802 527 825 547
rect 760 497 825 527
rect 345 476 410 497
rect 300 413 410 476
rect 440 471 496 497
rect 440 437 451 471
rect 485 437 496 471
rect 440 413 496 437
rect 526 471 636 497
rect 526 437 589 471
rect 623 437 636 471
rect 526 413 636 437
rect 666 413 708 497
rect 738 413 825 497
rect 760 379 825 413
rect 855 421 927 547
rect 855 387 866 421
rect 900 387 927 421
rect 855 379 927 387
rect 957 535 1064 547
rect 957 501 1022 535
rect 1056 501 1064 535
rect 957 463 1064 501
rect 1210 539 1267 547
rect 1210 505 1222 539
rect 1256 505 1267 539
rect 1210 463 1267 505
rect 957 425 1086 463
rect 957 391 1022 425
rect 1056 391 1086 425
rect 957 379 1086 391
rect 1116 379 1158 463
rect 1188 452 1267 463
rect 1188 418 1223 452
rect 1257 418 1267 452
rect 1188 379 1267 418
rect 1297 534 1350 547
rect 1297 500 1308 534
rect 1342 500 1350 534
rect 1297 425 1350 500
rect 1297 391 1308 425
rect 1342 391 1350 425
rect 1297 379 1350 391
rect 1469 512 1522 573
rect 1469 478 1477 512
rect 1511 478 1522 512
rect 1469 415 1522 478
rect 1469 381 1477 415
rect 1511 381 1522 415
rect 1469 367 1522 381
rect 1552 599 1605 619
rect 1552 565 1563 599
rect 1597 565 1605 599
rect 1552 502 1605 565
rect 1552 468 1563 502
rect 1597 468 1605 502
rect 1552 420 1605 468
rect 1552 386 1563 420
rect 1597 386 1605 420
rect 1552 367 1605 386
<< ndiffc >>
rect 248 187 282 221
rect 358 171 392 205
rect 465 188 499 222
rect 551 188 585 222
rect 35 95 69 129
rect 121 96 155 130
rect 730 148 764 182
rect 798 148 832 182
rect 891 199 925 233
rect 897 131 931 165
rect 1014 144 1048 178
rect 1211 155 1245 189
rect 1211 87 1245 121
rect 1311 155 1345 189
rect 1311 87 1345 121
rect 1477 169 1511 203
rect 1477 59 1511 93
rect 1563 169 1597 203
rect 1563 67 1597 101
<< pdiffc >>
rect 35 550 69 584
rect 35 481 69 515
rect 121 548 155 582
rect 121 480 155 514
rect 225 493 259 527
rect 225 425 259 459
rect 311 476 345 510
rect 768 527 802 561
rect 1477 573 1511 607
rect 451 437 485 471
rect 589 437 623 471
rect 866 387 900 421
rect 1022 501 1056 535
rect 1222 505 1256 539
rect 1022 391 1056 425
rect 1223 418 1257 452
rect 1308 500 1342 534
rect 1308 391 1342 425
rect 1477 478 1511 512
rect 1477 381 1511 415
rect 1563 565 1597 599
rect 1563 468 1597 502
rect 1563 386 1597 420
<< poly >>
rect 80 596 110 622
rect 270 615 957 645
rect 1522 619 1552 645
rect 270 541 300 615
rect 80 403 110 468
rect 410 497 440 523
rect 496 497 526 523
rect 636 497 666 615
rect 825 547 855 573
rect 927 547 957 615
rect 1107 586 1188 602
rect 1107 552 1126 586
rect 1160 552 1188 586
rect 708 497 738 523
rect 67 373 110 403
rect 67 325 97 373
rect 270 325 300 413
rect 410 335 440 413
rect 496 381 526 413
rect 636 387 666 413
rect 496 365 571 381
rect 31 309 110 325
rect 31 275 47 309
rect 81 275 110 309
rect 31 241 110 275
rect 31 207 47 241
rect 81 207 110 241
rect 31 191 110 207
rect 152 309 323 325
rect 152 275 168 309
rect 202 295 323 309
rect 202 275 218 295
rect 152 241 218 275
rect 293 247 323 295
rect 365 319 454 335
rect 365 285 381 319
rect 415 285 454 319
rect 496 331 521 365
rect 555 345 571 365
rect 555 331 626 345
rect 708 339 738 413
rect 1107 536 1188 552
rect 1267 547 1297 573
rect 1086 463 1116 489
rect 1158 463 1188 536
rect 496 315 626 331
rect 365 269 454 285
rect 424 247 454 269
rect 510 247 540 273
rect 596 247 626 315
rect 674 323 740 339
rect 825 335 855 379
rect 927 353 957 379
rect 674 303 690 323
rect 668 289 690 303
rect 724 289 740 323
rect 668 273 740 289
rect 796 319 880 335
rect 796 285 812 319
rect 846 285 880 319
rect 1086 307 1116 379
rect 1005 305 1116 307
rect 668 247 698 273
rect 796 269 880 285
rect 850 247 880 269
rect 948 289 1116 305
rect 948 255 971 289
rect 1005 277 1116 289
rect 1005 255 1035 277
rect 152 207 168 241
rect 202 207 218 241
rect 152 191 218 207
rect 80 154 110 191
rect 80 44 110 70
rect 293 51 323 163
rect 424 137 454 163
rect 510 51 540 163
rect 596 137 626 163
rect 668 137 698 163
rect 948 239 1035 255
rect 948 203 978 239
rect 1086 203 1116 229
rect 1158 203 1188 379
rect 1267 294 1297 379
rect 1522 331 1552 367
rect 1459 304 1552 331
rect 1245 291 1317 294
rect 1245 277 1319 291
rect 1245 242 1263 277
rect 1299 242 1319 277
rect 1459 270 1487 304
rect 1521 270 1552 304
rect 1459 250 1552 270
rect 1245 224 1319 242
rect 1259 203 1289 224
rect 1522 215 1552 250
rect 850 93 880 119
rect 948 93 978 119
rect 1086 51 1116 119
rect 1158 93 1188 119
rect 293 21 1116 51
rect 1259 49 1289 75
rect 1522 21 1552 47
<< polycont >>
rect 1126 552 1160 586
rect 47 275 81 309
rect 47 207 81 241
rect 168 275 202 309
rect 381 285 415 319
rect 521 331 555 365
rect 690 289 724 323
rect 812 285 846 319
rect 971 255 1005 289
rect 168 207 202 241
rect 1263 242 1299 277
rect 1487 270 1521 304
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 584 85 649
rect 19 550 35 584
rect 69 550 85 584
rect 19 515 85 550
rect 19 481 35 515
rect 69 481 85 515
rect 19 465 85 481
rect 119 582 159 598
rect 119 548 121 582
rect 155 548 159 582
rect 119 514 159 548
rect 119 480 121 514
rect 155 480 159 514
rect 17 309 85 431
rect 17 275 47 309
rect 81 275 85 309
rect 17 241 85 275
rect 17 207 47 241
rect 81 207 85 241
rect 17 168 85 207
rect 119 325 159 480
rect 209 527 270 543
rect 209 493 225 527
rect 259 493 270 527
rect 209 459 270 493
rect 304 510 347 649
rect 304 476 311 510
rect 345 476 347 510
rect 304 460 347 476
rect 381 521 699 576
rect 752 561 818 649
rect 752 527 768 561
rect 802 527 818 561
rect 1110 586 1177 597
rect 1110 552 1126 586
rect 1160 552 1177 586
rect 1022 535 1075 551
rect 1110 541 1177 552
rect 209 425 225 459
rect 259 426 270 459
rect 381 426 415 521
rect 259 425 415 426
rect 209 409 415 425
rect 236 392 415 409
rect 449 471 485 487
rect 449 437 451 471
rect 119 309 202 325
rect 119 275 168 309
rect 119 241 202 275
rect 119 207 168 241
rect 119 191 202 207
rect 236 221 282 392
rect 325 319 415 358
rect 325 285 381 319
rect 325 242 415 285
rect 19 129 85 134
rect 19 95 35 129
rect 69 95 85 129
rect 19 17 85 95
rect 119 130 171 191
rect 236 187 248 221
rect 449 238 485 437
rect 519 365 555 521
rect 665 491 699 521
rect 1056 501 1075 535
rect 519 331 521 365
rect 519 315 555 331
rect 589 471 631 487
rect 623 437 631 471
rect 665 457 986 491
rect 589 255 631 437
rect 674 421 916 423
rect 674 387 866 421
rect 900 387 916 421
rect 674 371 916 387
rect 674 323 740 371
rect 674 289 690 323
rect 724 289 740 323
rect 796 319 848 335
rect 796 285 812 319
rect 846 285 848 319
rect 796 255 848 285
rect 589 238 848 255
rect 449 222 515 238
rect 236 171 282 187
rect 342 205 408 208
rect 342 171 358 205
rect 392 171 408 205
rect 449 188 465 222
rect 499 188 515 222
rect 449 172 515 188
rect 551 222 848 238
rect 585 221 848 222
rect 882 249 916 371
rect 952 319 986 457
rect 1022 425 1075 501
rect 1056 391 1075 425
rect 1022 375 1075 391
rect 952 289 1007 319
rect 952 285 971 289
rect 1005 255 1007 289
rect 882 233 937 249
rect 971 239 1007 255
rect 1041 259 1075 375
rect 1135 359 1170 541
rect 1212 539 1272 649
rect 1461 607 1521 649
rect 1461 573 1477 607
rect 1511 573 1521 607
rect 1212 505 1222 539
rect 1256 505 1272 539
rect 1212 452 1272 505
rect 1212 418 1223 452
rect 1257 418 1272 452
rect 1212 393 1272 418
rect 1308 534 1397 550
rect 1342 500 1397 534
rect 1308 425 1397 500
rect 1342 391 1397 425
rect 1308 359 1397 391
rect 1461 512 1521 573
rect 1461 478 1477 512
rect 1511 478 1521 512
rect 1461 415 1521 478
rect 1461 381 1477 415
rect 1511 381 1521 415
rect 1461 365 1521 381
rect 1555 599 1613 615
rect 1555 565 1563 599
rect 1597 565 1613 599
rect 1555 502 1613 565
rect 1555 468 1563 502
rect 1597 468 1613 502
rect 1555 420 1613 468
rect 1555 386 1563 420
rect 1597 386 1613 420
rect 1135 331 1397 359
rect 1135 325 1521 331
rect 1363 304 1521 325
rect 1245 277 1319 291
rect 1245 259 1263 277
rect 1041 242 1263 259
rect 1299 242 1319 277
rect 585 188 625 221
rect 551 172 625 188
rect 882 199 891 233
rect 925 199 937 233
rect 714 182 848 187
rect 119 96 121 130
rect 155 96 171 130
rect 119 80 171 96
rect 342 17 408 171
rect 714 148 730 182
rect 764 148 798 182
rect 832 148 848 182
rect 714 17 848 148
rect 882 165 937 199
rect 1041 225 1319 242
rect 1041 194 1079 225
rect 1245 224 1319 225
rect 1363 270 1487 304
rect 1363 254 1521 270
rect 882 131 897 165
rect 931 131 937 165
rect 882 115 937 131
rect 998 178 1079 194
rect 1363 189 1434 254
rect 998 144 1014 178
rect 1048 144 1079 178
rect 998 128 1079 144
rect 1195 155 1211 189
rect 1245 155 1261 189
rect 1195 121 1261 155
rect 1195 87 1211 121
rect 1245 87 1261 121
rect 1195 17 1261 87
rect 1295 155 1311 189
rect 1345 155 1434 189
rect 1295 121 1434 155
rect 1295 87 1311 121
rect 1345 87 1434 121
rect 1295 83 1434 87
rect 1468 203 1521 219
rect 1468 169 1477 203
rect 1511 169 1521 203
rect 1468 93 1521 169
rect 1468 59 1477 93
rect 1511 59 1521 93
rect 1468 17 1521 59
rect 1555 203 1613 386
rect 1555 169 1563 203
rect 1597 169 1613 203
rect 1555 101 1613 169
rect 1555 67 1563 101
rect 1597 67 1613 101
rect 1555 51 1613 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxtp_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFclass CORE
string LEFsite unit
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string GDS_START 110132
string GDS_END 122576
string LEFsymmetry X Y R90
<< end >>
