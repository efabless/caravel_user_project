magic
tech sky130A
magscale 1 2
timestamp 1619036415
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 106 484 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10230 119200 10286 120000
rect 11794 119200 11850 120000
rect 13358 119200 13414 120000
rect 14922 119200 14978 120000
rect 16486 119200 16542 120000
rect 18050 119200 18106 120000
rect 19706 119200 19762 120000
rect 21270 119200 21326 120000
rect 22834 119200 22890 120000
rect 24398 119200 24454 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 29182 119200 29238 120000
rect 30746 119200 30802 120000
rect 32310 119200 32366 120000
rect 33874 119200 33930 120000
rect 35438 119200 35494 120000
rect 37002 119200 37058 120000
rect 38658 119200 38714 120000
rect 40222 119200 40278 120000
rect 41786 119200 41842 120000
rect 43350 119200 43406 120000
rect 44914 119200 44970 120000
rect 46478 119200 46534 120000
rect 48134 119200 48190 120000
rect 49698 119200 49754 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54390 119200 54446 120000
rect 55954 119200 56010 120000
rect 57610 119200 57666 120000
rect 59174 119200 59230 120000
rect 60738 119200 60794 120000
rect 62302 119200 62358 120000
rect 63866 119200 63922 120000
rect 65430 119200 65486 120000
rect 67086 119200 67142 120000
rect 68650 119200 68706 120000
rect 70214 119200 70270 120000
rect 71778 119200 71834 120000
rect 73342 119200 73398 120000
rect 74906 119200 74962 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79690 119200 79746 120000
rect 81254 119200 81310 120000
rect 82818 119200 82874 120000
rect 84382 119200 84438 120000
rect 86038 119200 86094 120000
rect 87602 119200 87658 120000
rect 89166 119200 89222 120000
rect 90730 119200 90786 120000
rect 92294 119200 92350 120000
rect 93858 119200 93914 120000
rect 95514 119200 95570 120000
rect 97078 119200 97134 120000
rect 98642 119200 98698 120000
rect 100206 119200 100262 120000
rect 101770 119200 101826 120000
rect 103334 119200 103390 120000
rect 104990 119200 105046 120000
rect 106554 119200 106610 120000
rect 108118 119200 108174 120000
rect 109682 119200 109738 120000
rect 111246 119200 111302 120000
rect 112810 119200 112866 120000
rect 114466 119200 114522 120000
rect 116030 119200 116086 120000
rect 117594 119200 117650 120000
rect 119158 119200 119214 120000
rect 120722 119200 120778 120000
rect 122286 119200 122342 120000
rect 123942 119200 123998 120000
rect 125506 119200 125562 120000
rect 127070 119200 127126 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131762 119200 131818 120000
rect 133418 119200 133474 120000
rect 134982 119200 135038 120000
rect 136546 119200 136602 120000
rect 138110 119200 138166 120000
rect 139674 119200 139730 120000
rect 141238 119200 141294 120000
rect 142894 119200 142950 120000
rect 144458 119200 144514 120000
rect 146022 119200 146078 120000
rect 147586 119200 147642 120000
rect 149150 119200 149206 120000
rect 150714 119200 150770 120000
rect 152370 119200 152426 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 157062 119200 157118 120000
rect 158626 119200 158682 120000
rect 160190 119200 160246 120000
rect 161846 119200 161902 120000
rect 163410 119200 163466 120000
rect 164974 119200 165030 120000
rect 166538 119200 166594 120000
rect 168102 119200 168158 120000
rect 169666 119200 169722 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119200
rect 866 119144 2262 119200
rect 2430 119144 3826 119200
rect 3994 119144 5390 119200
rect 5558 119144 6954 119200
rect 7122 119144 8518 119200
rect 8686 119144 10174 119200
rect 10342 119144 11738 119200
rect 11906 119144 13302 119200
rect 13470 119144 14866 119200
rect 15034 119144 16430 119200
rect 16598 119144 17994 119200
rect 18162 119144 19650 119200
rect 19818 119144 21214 119200
rect 21382 119144 22778 119200
rect 22946 119144 24342 119200
rect 24510 119144 25906 119200
rect 26074 119144 27470 119200
rect 27638 119144 29126 119200
rect 29294 119144 30690 119200
rect 30858 119144 32254 119200
rect 32422 119144 33818 119200
rect 33986 119144 35382 119200
rect 35550 119144 36946 119200
rect 37114 119144 38602 119200
rect 38770 119144 40166 119200
rect 40334 119144 41730 119200
rect 41898 119144 43294 119200
rect 43462 119144 44858 119200
rect 45026 119144 46422 119200
rect 46590 119144 48078 119200
rect 48246 119144 49642 119200
rect 49810 119144 51206 119200
rect 51374 119144 52770 119200
rect 52938 119144 54334 119200
rect 54502 119144 55898 119200
rect 56066 119144 57554 119200
rect 57722 119144 59118 119200
rect 59286 119144 60682 119200
rect 60850 119144 62246 119200
rect 62414 119144 63810 119200
rect 63978 119144 65374 119200
rect 65542 119144 67030 119200
rect 67198 119144 68594 119200
rect 68762 119144 70158 119200
rect 70326 119144 71722 119200
rect 71890 119144 73286 119200
rect 73454 119144 74850 119200
rect 75018 119144 76506 119200
rect 76674 119144 78070 119200
rect 78238 119144 79634 119200
rect 79802 119144 81198 119200
rect 81366 119144 82762 119200
rect 82930 119144 84326 119200
rect 84494 119144 85982 119200
rect 86150 119144 87546 119200
rect 87714 119144 89110 119200
rect 89278 119144 90674 119200
rect 90842 119144 92238 119200
rect 92406 119144 93802 119200
rect 93970 119144 95458 119200
rect 95626 119144 97022 119200
rect 97190 119144 98586 119200
rect 98754 119144 100150 119200
rect 100318 119144 101714 119200
rect 101882 119144 103278 119200
rect 103446 119144 104934 119200
rect 105102 119144 106498 119200
rect 106666 119144 108062 119200
rect 108230 119144 109626 119200
rect 109794 119144 111190 119200
rect 111358 119144 112754 119200
rect 112922 119144 114410 119200
rect 114578 119144 115974 119200
rect 116142 119144 117538 119200
rect 117706 119144 119102 119200
rect 119270 119144 120666 119200
rect 120834 119144 122230 119200
rect 122398 119144 123886 119200
rect 124054 119144 125450 119200
rect 125618 119144 127014 119200
rect 127182 119144 128578 119200
rect 128746 119144 130142 119200
rect 130310 119144 131706 119200
rect 131874 119144 133362 119200
rect 133530 119144 134926 119200
rect 135094 119144 136490 119200
rect 136658 119144 138054 119200
rect 138222 119144 139618 119200
rect 139786 119144 141182 119200
rect 141350 119144 142838 119200
rect 143006 119144 144402 119200
rect 144570 119144 145966 119200
rect 146134 119144 147530 119200
rect 147698 119144 149094 119200
rect 149262 119144 150658 119200
rect 150826 119144 152314 119200
rect 152482 119144 153878 119200
rect 154046 119144 155442 119200
rect 155610 119144 157006 119200
rect 157174 119144 158570 119200
rect 158738 119144 160134 119200
rect 160302 119144 161790 119200
rect 161958 119144 163354 119200
rect 163522 119144 164918 119200
rect 165086 119144 166482 119200
rect 166650 119144 168046 119200
rect 168214 119144 169610 119200
rect 169778 119144 171266 119200
rect 171434 119144 172830 119200
rect 172998 119144 174394 119200
rect 174562 119144 175958 119200
rect 176126 119144 177522 119200
rect 177690 119144 179086 119200
rect 179254 119144 179840 119200
rect 112 856 179840 119144
rect 222 478 330 856
rect 498 478 698 856
rect 866 478 1066 856
rect 1234 478 1434 856
rect 1602 478 1802 856
rect 1970 478 2170 856
rect 2338 478 2538 856
rect 2706 478 2906 856
rect 3074 478 3274 856
rect 3442 478 3642 856
rect 3810 478 4010 856
rect 4178 478 4378 856
rect 4546 478 4746 856
rect 4914 478 5114 856
rect 5282 478 5482 856
rect 5650 478 5850 856
rect 6018 478 6218 856
rect 6386 478 6586 856
rect 6754 478 6954 856
rect 7122 478 7322 856
rect 7490 478 7690 856
rect 7858 478 8058 856
rect 8226 478 8426 856
rect 8594 478 8794 856
rect 8962 478 9162 856
rect 9330 478 9530 856
rect 9698 478 9898 856
rect 10066 478 10266 856
rect 10434 478 10634 856
rect 10802 478 11002 856
rect 11170 478 11370 856
rect 11538 478 11738 856
rect 11906 478 12106 856
rect 12274 478 12474 856
rect 12642 478 12842 856
rect 13010 478 13210 856
rect 13378 478 13578 856
rect 13746 478 13946 856
rect 14114 478 14314 856
rect 14482 478 14682 856
rect 14850 478 15050 856
rect 15218 478 15418 856
rect 15586 478 15786 856
rect 15954 478 16154 856
rect 16322 478 16522 856
rect 16690 478 16890 856
rect 17058 478 17258 856
rect 17426 478 17626 856
rect 17794 478 17994 856
rect 18162 478 18362 856
rect 18530 478 18730 856
rect 18898 478 19098 856
rect 19266 478 19466 856
rect 19634 478 19834 856
rect 20002 478 20202 856
rect 20370 478 20570 856
rect 20738 478 20938 856
rect 21106 478 21306 856
rect 21474 478 21674 856
rect 21842 478 22042 856
rect 22210 478 22410 856
rect 22578 478 22778 856
rect 22946 478 23146 856
rect 23314 478 23514 856
rect 23682 478 23882 856
rect 24050 478 24250 856
rect 24418 478 24618 856
rect 24786 478 24986 856
rect 25154 478 25354 856
rect 25522 478 25722 856
rect 25890 478 26090 856
rect 26258 478 26458 856
rect 26626 478 26826 856
rect 26994 478 27194 856
rect 27362 478 27562 856
rect 27730 478 27930 856
rect 28098 478 28298 856
rect 28466 478 28666 856
rect 28834 478 29034 856
rect 29202 478 29402 856
rect 29570 478 29770 856
rect 29938 478 30138 856
rect 30306 478 30506 856
rect 30674 478 30874 856
rect 31042 478 31242 856
rect 31410 478 31610 856
rect 31778 478 31978 856
rect 32146 478 32346 856
rect 32514 478 32714 856
rect 32882 478 33082 856
rect 33250 478 33450 856
rect 33618 478 33818 856
rect 33986 478 34186 856
rect 34354 478 34554 856
rect 34722 478 34922 856
rect 35090 478 35290 856
rect 35458 478 35658 856
rect 35826 478 36026 856
rect 36194 478 36394 856
rect 36562 478 36762 856
rect 36930 478 37130 856
rect 37298 478 37498 856
rect 37666 478 37866 856
rect 38034 478 38234 856
rect 38402 478 38602 856
rect 38770 478 38970 856
rect 39138 478 39338 856
rect 39506 478 39706 856
rect 39874 478 40074 856
rect 40242 478 40442 856
rect 40610 478 40810 856
rect 40978 478 41178 856
rect 41346 478 41546 856
rect 41714 478 41914 856
rect 42082 478 42282 856
rect 42450 478 42650 856
rect 42818 478 43018 856
rect 43186 478 43386 856
rect 43554 478 43754 856
rect 43922 478 44122 856
rect 44290 478 44490 856
rect 44658 478 44858 856
rect 45026 478 45226 856
rect 45394 478 45594 856
rect 45762 478 45962 856
rect 46130 478 46330 856
rect 46498 478 46698 856
rect 46866 478 47066 856
rect 47234 478 47434 856
rect 47602 478 47802 856
rect 47970 478 48170 856
rect 48338 478 48538 856
rect 48706 478 48906 856
rect 49074 478 49274 856
rect 49442 478 49642 856
rect 49810 478 50010 856
rect 50178 478 50378 856
rect 50546 478 50746 856
rect 50914 478 51114 856
rect 51282 478 51482 856
rect 51650 478 51850 856
rect 52018 478 52218 856
rect 52386 478 52586 856
rect 52754 478 52954 856
rect 53122 478 53322 856
rect 53490 478 53690 856
rect 53858 478 54058 856
rect 54226 478 54426 856
rect 54594 478 54794 856
rect 54962 478 55162 856
rect 55330 478 55530 856
rect 55698 478 55898 856
rect 56066 478 56266 856
rect 56434 478 56634 856
rect 56802 478 57002 856
rect 57170 478 57370 856
rect 57538 478 57738 856
rect 57906 478 58106 856
rect 58274 478 58474 856
rect 58642 478 58842 856
rect 59010 478 59210 856
rect 59378 478 59578 856
rect 59746 478 59946 856
rect 60114 478 60222 856
rect 60390 478 60590 856
rect 60758 478 60958 856
rect 61126 478 61326 856
rect 61494 478 61694 856
rect 61862 478 62062 856
rect 62230 478 62430 856
rect 62598 478 62798 856
rect 62966 478 63166 856
rect 63334 478 63534 856
rect 63702 478 63902 856
rect 64070 478 64270 856
rect 64438 478 64638 856
rect 64806 478 65006 856
rect 65174 478 65374 856
rect 65542 478 65742 856
rect 65910 478 66110 856
rect 66278 478 66478 856
rect 66646 478 66846 856
rect 67014 478 67214 856
rect 67382 478 67582 856
rect 67750 478 67950 856
rect 68118 478 68318 856
rect 68486 478 68686 856
rect 68854 478 69054 856
rect 69222 478 69422 856
rect 69590 478 69790 856
rect 69958 478 70158 856
rect 70326 478 70526 856
rect 70694 478 70894 856
rect 71062 478 71262 856
rect 71430 478 71630 856
rect 71798 478 71998 856
rect 72166 478 72366 856
rect 72534 478 72734 856
rect 72902 478 73102 856
rect 73270 478 73470 856
rect 73638 478 73838 856
rect 74006 478 74206 856
rect 74374 478 74574 856
rect 74742 478 74942 856
rect 75110 478 75310 856
rect 75478 478 75678 856
rect 75846 478 76046 856
rect 76214 478 76414 856
rect 76582 478 76782 856
rect 76950 478 77150 856
rect 77318 478 77518 856
rect 77686 478 77886 856
rect 78054 478 78254 856
rect 78422 478 78622 856
rect 78790 478 78990 856
rect 79158 478 79358 856
rect 79526 478 79726 856
rect 79894 478 80094 856
rect 80262 478 80462 856
rect 80630 478 80830 856
rect 80998 478 81198 856
rect 81366 478 81566 856
rect 81734 478 81934 856
rect 82102 478 82302 856
rect 82470 478 82670 856
rect 82838 478 83038 856
rect 83206 478 83406 856
rect 83574 478 83774 856
rect 83942 478 84142 856
rect 84310 478 84510 856
rect 84678 478 84878 856
rect 85046 478 85246 856
rect 85414 478 85614 856
rect 85782 478 85982 856
rect 86150 478 86350 856
rect 86518 478 86718 856
rect 86886 478 87086 856
rect 87254 478 87454 856
rect 87622 478 87822 856
rect 87990 478 88190 856
rect 88358 478 88558 856
rect 88726 478 88926 856
rect 89094 478 89294 856
rect 89462 478 89662 856
rect 89830 478 90030 856
rect 90198 478 90398 856
rect 90566 478 90766 856
rect 90934 478 91134 856
rect 91302 478 91502 856
rect 91670 478 91870 856
rect 92038 478 92238 856
rect 92406 478 92606 856
rect 92774 478 92974 856
rect 93142 478 93342 856
rect 93510 478 93710 856
rect 93878 478 94078 856
rect 94246 478 94446 856
rect 94614 478 94814 856
rect 94982 478 95182 856
rect 95350 478 95550 856
rect 95718 478 95918 856
rect 96086 478 96286 856
rect 96454 478 96654 856
rect 96822 478 97022 856
rect 97190 478 97390 856
rect 97558 478 97758 856
rect 97926 478 98126 856
rect 98294 478 98494 856
rect 98662 478 98862 856
rect 99030 478 99230 856
rect 99398 478 99598 856
rect 99766 478 99966 856
rect 100134 478 100334 856
rect 100502 478 100702 856
rect 100870 478 101070 856
rect 101238 478 101438 856
rect 101606 478 101806 856
rect 101974 478 102174 856
rect 102342 478 102542 856
rect 102710 478 102910 856
rect 103078 478 103278 856
rect 103446 478 103646 856
rect 103814 478 104014 856
rect 104182 478 104382 856
rect 104550 478 104750 856
rect 104918 478 105118 856
rect 105286 478 105486 856
rect 105654 478 105854 856
rect 106022 478 106222 856
rect 106390 478 106590 856
rect 106758 478 106958 856
rect 107126 478 107326 856
rect 107494 478 107694 856
rect 107862 478 108062 856
rect 108230 478 108430 856
rect 108598 478 108798 856
rect 108966 478 109166 856
rect 109334 478 109534 856
rect 109702 478 109902 856
rect 110070 478 110270 856
rect 110438 478 110638 856
rect 110806 478 111006 856
rect 111174 478 111374 856
rect 111542 478 111742 856
rect 111910 478 112110 856
rect 112278 478 112478 856
rect 112646 478 112846 856
rect 113014 478 113214 856
rect 113382 478 113582 856
rect 113750 478 113950 856
rect 114118 478 114318 856
rect 114486 478 114686 856
rect 114854 478 115054 856
rect 115222 478 115422 856
rect 115590 478 115790 856
rect 115958 478 116158 856
rect 116326 478 116526 856
rect 116694 478 116894 856
rect 117062 478 117262 856
rect 117430 478 117630 856
rect 117798 478 117998 856
rect 118166 478 118366 856
rect 118534 478 118734 856
rect 118902 478 119102 856
rect 119270 478 119470 856
rect 119638 478 119838 856
rect 120006 478 120114 856
rect 120282 478 120482 856
rect 120650 478 120850 856
rect 121018 478 121218 856
rect 121386 478 121586 856
rect 121754 478 121954 856
rect 122122 478 122322 856
rect 122490 478 122690 856
rect 122858 478 123058 856
rect 123226 478 123426 856
rect 123594 478 123794 856
rect 123962 478 124162 856
rect 124330 478 124530 856
rect 124698 478 124898 856
rect 125066 478 125266 856
rect 125434 478 125634 856
rect 125802 478 126002 856
rect 126170 478 126370 856
rect 126538 478 126738 856
rect 126906 478 127106 856
rect 127274 478 127474 856
rect 127642 478 127842 856
rect 128010 478 128210 856
rect 128378 478 128578 856
rect 128746 478 128946 856
rect 129114 478 129314 856
rect 129482 478 129682 856
rect 129850 478 130050 856
rect 130218 478 130418 856
rect 130586 478 130786 856
rect 130954 478 131154 856
rect 131322 478 131522 856
rect 131690 478 131890 856
rect 132058 478 132258 856
rect 132426 478 132626 856
rect 132794 478 132994 856
rect 133162 478 133362 856
rect 133530 478 133730 856
rect 133898 478 134098 856
rect 134266 478 134466 856
rect 134634 478 134834 856
rect 135002 478 135202 856
rect 135370 478 135570 856
rect 135738 478 135938 856
rect 136106 478 136306 856
rect 136474 478 136674 856
rect 136842 478 137042 856
rect 137210 478 137410 856
rect 137578 478 137778 856
rect 137946 478 138146 856
rect 138314 478 138514 856
rect 138682 478 138882 856
rect 139050 478 139250 856
rect 139418 478 139618 856
rect 139786 478 139986 856
rect 140154 478 140354 856
rect 140522 478 140722 856
rect 140890 478 141090 856
rect 141258 478 141458 856
rect 141626 478 141826 856
rect 141994 478 142194 856
rect 142362 478 142562 856
rect 142730 478 142930 856
rect 143098 478 143298 856
rect 143466 478 143666 856
rect 143834 478 144034 856
rect 144202 478 144402 856
rect 144570 478 144770 856
rect 144938 478 145138 856
rect 145306 478 145506 856
rect 145674 478 145874 856
rect 146042 478 146242 856
rect 146410 478 146610 856
rect 146778 478 146978 856
rect 147146 478 147346 856
rect 147514 478 147714 856
rect 147882 478 148082 856
rect 148250 478 148450 856
rect 148618 478 148818 856
rect 148986 478 149186 856
rect 149354 478 149554 856
rect 149722 478 149922 856
rect 150090 478 150290 856
rect 150458 478 150658 856
rect 150826 478 151026 856
rect 151194 478 151394 856
rect 151562 478 151762 856
rect 151930 478 152130 856
rect 152298 478 152498 856
rect 152666 478 152866 856
rect 153034 478 153234 856
rect 153402 478 153602 856
rect 153770 478 153970 856
rect 154138 478 154338 856
rect 154506 478 154706 856
rect 154874 478 155074 856
rect 155242 478 155442 856
rect 155610 478 155810 856
rect 155978 478 156178 856
rect 156346 478 156546 856
rect 156714 478 156914 856
rect 157082 478 157282 856
rect 157450 478 157650 856
rect 157818 478 158018 856
rect 158186 478 158386 856
rect 158554 478 158754 856
rect 158922 478 159122 856
rect 159290 478 159490 856
rect 159658 478 159858 856
rect 160026 478 160226 856
rect 160394 478 160594 856
rect 160762 478 160962 856
rect 161130 478 161330 856
rect 161498 478 161698 856
rect 161866 478 162066 856
rect 162234 478 162434 856
rect 162602 478 162802 856
rect 162970 478 163170 856
rect 163338 478 163538 856
rect 163706 478 163906 856
rect 164074 478 164274 856
rect 164442 478 164642 856
rect 164810 478 165010 856
rect 165178 478 165378 856
rect 165546 478 165746 856
rect 165914 478 166114 856
rect 166282 478 166482 856
rect 166650 478 166850 856
rect 167018 478 167218 856
rect 167386 478 167586 856
rect 167754 478 167954 856
rect 168122 478 168322 856
rect 168490 478 168690 856
rect 168858 478 169058 856
rect 169226 478 169426 856
rect 169594 478 169794 856
rect 169962 478 170162 856
rect 170330 478 170530 856
rect 170698 478 170898 856
rect 171066 478 171266 856
rect 171434 478 171634 856
rect 171802 478 172002 856
rect 172170 478 172370 856
rect 172538 478 172738 856
rect 172906 478 173106 856
rect 173274 478 173474 856
rect 173642 478 173842 856
rect 174010 478 174210 856
rect 174378 478 174578 856
rect 174746 478 174946 856
rect 175114 478 175314 856
rect 175482 478 175682 856
rect 175850 478 176050 856
rect 176218 478 176418 856
rect 176586 478 176786 856
rect 176954 478 177154 856
rect 177322 478 177522 856
rect 177690 478 177890 856
rect 178058 478 178258 856
rect 178426 478 178626 856
rect 178794 478 178994 856
rect 179162 478 179362 856
rect 179530 478 179730 856
<< obsm3 >>
rect 1669 1803 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 2550 2048 4128 5541
rect 4608 2096 4788 5541
rect 5268 2096 5448 5541
rect 5928 2096 6108 5541
rect 6588 2096 19488 5541
rect 4608 2048 19488 2096
rect 19968 2096 20148 5541
rect 20628 2096 20808 5541
rect 21288 2096 21468 5541
rect 21948 2096 34848 5541
rect 19968 2048 34848 2096
rect 35328 2096 35508 5541
rect 35988 2096 36168 5541
rect 36648 2096 36828 5541
rect 37308 2096 50208 5541
rect 35328 2048 50208 2096
rect 50688 2096 50868 5541
rect 51348 2096 51528 5541
rect 52008 2096 52188 5541
rect 52668 2096 65568 5541
rect 50688 2048 65568 2096
rect 66048 2096 66228 5541
rect 66708 2096 66888 5541
rect 67368 2096 67548 5541
rect 68028 2096 80928 5541
rect 66048 2048 80928 2096
rect 81408 2096 81588 5541
rect 82068 2096 82248 5541
rect 82728 2096 82908 5541
rect 83388 2096 96288 5541
rect 81408 2048 96288 2096
rect 96768 2096 96948 5541
rect 97428 2096 97608 5541
rect 98088 2096 98268 5541
rect 98748 2096 102330 5541
rect 96768 2048 102330 2096
rect 2550 1803 102330 2048
<< obsm5 >>
rect 2508 2900 102372 3220
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 48134 119200 48190 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52826 119200 52882 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57610 119200 57666 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 62302 119200 62358 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 67086 119200 67142 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71778 119200 71834 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 81254 119200 81310 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 95514 119200 95570 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 100206 119200 100262 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104990 119200 105046 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 109682 119200 109738 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 114466 119200 114522 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 123942 119200 123998 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 128634 119200 128690 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 133418 119200 133474 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 138110 119200 138166 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10230 119200 10286 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 142894 119200 142950 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 147586 119200 147642 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 152370 119200 152426 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 157062 119200 157118 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 161846 119200 161902 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 166538 119200 166594 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 171322 119200 171378 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 176014 119200 176070 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14922 119200 14978 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19706 119200 19762 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24398 119200 24454 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 29182 119200 29238 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33874 119200 33930 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38658 119200 38714 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 43350 119200 43406 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49698 119200 49754 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 54390 119200 54446 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 59174 119200 59230 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63866 119200 63922 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 73342 119200 73398 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82818 119200 82874 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 92294 119200 92350 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 97078 119200 97134 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 111246 119200 111302 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 116030 119200 116086 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 120722 119200 120778 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 125506 119200 125562 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 130198 119200 130254 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 139674 119200 139730 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11794 119200 11850 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 144458 119200 144514 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 149150 119200 149206 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 158626 119200 158682 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 163410 119200 163466 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 168102 119200 168158 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 172886 119200 172942 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16486 119200 16542 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21270 119200 21326 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35438 119200 35494 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 40222 119200 40278 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44914 119200 44970 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55954 119200 56010 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 65430 119200 65486 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 70214 119200 70270 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74906 119200 74962 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 79690 119200 79746 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 98642 119200 98698 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 103334 119200 103390 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 108118 119200 108174 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 112810 119200 112866 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 117594 119200 117650 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 122286 119200 122342 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 127070 119200 127126 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 131762 119200 131818 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 136546 119200 136602 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 141238 119200 141294 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13358 119200 13414 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 146022 119200 146078 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 150714 119200 150770 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 160190 119200 160246 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 164974 119200 165030 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 169666 119200 169722 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 174450 119200 174506 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 179142 119200 179198 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 18050 119200 18106 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22834 119200 22890 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27526 119200 27582 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32310 119200 32366 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37002 119200 37058 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41786 119200 41842 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46478 119200 46534 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 95606 0 95662 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 499 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 500 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 501 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 502 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 503 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 504 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[12]
port 505 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[13]
port 506 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[14]
port 507 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[15]
port 508 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[16]
port 509 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[17]
port 510 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[18]
port 511 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[19]
port 512 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 513 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[20]
port 514 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[21]
port 515 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[22]
port 516 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[23]
port 517 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_adr_i[24]
port 518 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[25]
port 519 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[26]
port 520 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[27]
port 521 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[28]
port 522 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[29]
port 523 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 524 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_adr_i[30]
port 525 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[31]
port 526 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 527 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 528 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 529 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 530 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 531 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 532 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 533 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 534 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 535 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 536 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 537 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[12]
port 538 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[13]
port 539 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[14]
port 540 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[15]
port 541 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[16]
port 542 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[17]
port 543 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[18]
port 544 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[19]
port 545 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 546 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[20]
port 547 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[21]
port 548 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[22]
port 549 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[23]
port 550 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[24]
port 551 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[25]
port 552 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[26]
port 553 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[27]
port 554 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[28]
port 555 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[29]
port 556 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 557 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[30]
port 558 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[31]
port 559 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 560 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 561 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 562 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 563 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 564 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 565 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 566 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 567 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 568 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[11]
port 569 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[12]
port 570 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[13]
port 571 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[14]
port 572 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[15]
port 573 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[16]
port 574 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[17]
port 575 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[18]
port 576 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[19]
port 577 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 578 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[20]
port 579 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[21]
port 580 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[22]
port 581 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_o[23]
port 582 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[24]
port 583 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[25]
port 584 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[26]
port 585 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[27]
port 586 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[28]
port 587 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[29]
port 588 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 589 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[30]
port 590 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_o[31]
port 591 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 592 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 593 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 594 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 595 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 596 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 597 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 598 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 599 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 600 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 601 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 602 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 603 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 604 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 606 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 607 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 611 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 619 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 623 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 624 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 625 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 629 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 630 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 631 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 635 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 636 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 637 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 641 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 642 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 643 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 647 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 648 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 649 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 652 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 7195308
string GDS_START 339680
<< end >>

