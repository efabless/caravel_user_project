magic
tech sky130A
timestamp 1640305290
<< metal1 >>
rect 475 555 525 605
rect -105 265 -55 275
rect -105 235 -95 265
rect -65 235 -55 265
rect -105 225 -55 235
rect 1055 265 1105 275
rect 1055 235 1065 265
rect 1095 235 1105 265
rect 1055 225 1105 235
<< via1 >>
rect -95 235 -65 265
rect 1065 235 1095 265
<< metal2 >>
rect 475 595 525 605
rect 475 565 485 595
rect 515 565 525 595
rect 475 555 525 565
rect -105 265 -55 275
rect -105 235 -95 265
rect -65 235 -55 265
rect -105 225 -55 235
rect 1055 265 1105 275
rect 1055 235 1065 265
rect 1095 235 1105 265
rect 1055 225 1105 235
rect 475 -65 525 -55
rect 475 -95 485 -65
rect 515 -95 525 -65
rect 475 -105 525 -95
<< via2 >>
rect 485 565 515 595
rect -95 235 -65 265
rect 1065 235 1095 265
rect 485 -95 515 -65
<< metal3 >>
rect 475 600 525 605
rect 475 560 480 600
rect 520 560 525 600
rect 475 555 525 560
rect -105 270 -55 275
rect -105 230 -100 270
rect -60 230 -55 270
rect -105 225 -55 230
rect -14 86 1014 514
rect 1055 270 1105 275
rect 1055 230 1060 270
rect 1100 230 1105 270
rect 1055 225 1105 230
rect -273 -14 1014 86
rect 475 -60 525 -55
rect 475 -100 480 -60
rect 520 -100 525 -60
rect 475 -105 525 -100
<< via3 >>
rect 480 595 520 600
rect 480 565 485 595
rect 485 565 515 595
rect 515 565 520 595
rect 480 560 520 565
rect -100 265 -60 270
rect -100 235 -95 265
rect -95 235 -65 265
rect -65 235 -60 265
rect -100 230 -60 235
rect 1060 265 1100 270
rect 1060 235 1065 265
rect 1065 235 1095 265
rect 1095 235 1100 265
rect 1060 230 1100 235
rect 480 -65 520 -60
rect 480 -95 485 -65
rect 485 -95 515 -65
rect 515 -95 520 -65
rect 480 -100 520 -95
<< mimcap >>
rect 0 300 1000 500
rect 0 200 450 300
rect 550 200 1000 300
rect 0 0 1000 200
<< mimcapcontact >>
rect 450 200 550 300
<< metal4 >>
rect 450 600 550 625
rect 450 560 480 600
rect 520 560 550 600
rect 450 300 550 560
rect -125 270 450 300
rect -125 230 -100 270
rect -60 230 450 270
rect -125 200 450 230
rect 550 270 1125 300
rect 550 230 1060 270
rect 1100 230 1125 270
rect 550 200 1125 230
rect 450 -60 550 200
rect 450 -100 480 -60
rect 520 -100 550 -60
rect 450 -125 550 -100
<< end >>
