magic
tech sky130A
magscale 1 2
timestamp 1621850781
<< obsli1 >>
rect 1104 1853 178848 117521
<< obsm1 >>
rect 106 1368 179846 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3882 119200 3938 120000
rect 5446 119200 5502 120000
rect 7010 119200 7066 120000
rect 8574 119200 8630 120000
rect 10138 119200 10194 120000
rect 11702 119200 11758 120000
rect 13266 119200 13322 120000
rect 14830 119200 14886 120000
rect 16394 119200 16450 120000
rect 17958 119200 18014 120000
rect 19522 119200 19578 120000
rect 21086 119200 21142 120000
rect 22650 119200 22706 120000
rect 24214 119200 24270 120000
rect 25778 119200 25834 120000
rect 27342 119200 27398 120000
rect 28906 119200 28962 120000
rect 30470 119200 30526 120000
rect 32034 119200 32090 120000
rect 33598 119200 33654 120000
rect 35162 119200 35218 120000
rect 36726 119200 36782 120000
rect 38290 119200 38346 120000
rect 39854 119200 39910 120000
rect 41418 119200 41474 120000
rect 42982 119200 43038 120000
rect 44546 119200 44602 120000
rect 46110 119200 46166 120000
rect 47674 119200 47730 120000
rect 49238 119200 49294 120000
rect 50802 119200 50858 120000
rect 52366 119200 52422 120000
rect 53930 119200 53986 120000
rect 55494 119200 55550 120000
rect 57058 119200 57114 120000
rect 58622 119200 58678 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63314 119200 63370 120000
rect 64878 119200 64934 120000
rect 66442 119200 66498 120000
rect 68006 119200 68062 120000
rect 69570 119200 69626 120000
rect 71134 119200 71190 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75826 119200 75882 120000
rect 77390 119200 77446 120000
rect 78954 119200 79010 120000
rect 80518 119200 80574 120000
rect 82082 119200 82138 120000
rect 83646 119200 83702 120000
rect 85210 119200 85266 120000
rect 86774 119200 86830 120000
rect 88338 119200 88394 120000
rect 89902 119200 89958 120000
rect 91558 119200 91614 120000
rect 93122 119200 93178 120000
rect 94686 119200 94742 120000
rect 96250 119200 96306 120000
rect 97814 119200 97870 120000
rect 99378 119200 99434 120000
rect 100942 119200 100998 120000
rect 102506 119200 102562 120000
rect 104070 119200 104126 120000
rect 105634 119200 105690 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110326 119200 110382 120000
rect 111890 119200 111946 120000
rect 113454 119200 113510 120000
rect 115018 119200 115074 120000
rect 116582 119200 116638 120000
rect 118146 119200 118202 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122838 119200 122894 120000
rect 124402 119200 124458 120000
rect 125966 119200 126022 120000
rect 127530 119200 127586 120000
rect 129094 119200 129150 120000
rect 130658 119200 130714 120000
rect 132222 119200 132278 120000
rect 133786 119200 133842 120000
rect 135350 119200 135406 120000
rect 136914 119200 136970 120000
rect 138478 119200 138534 120000
rect 140042 119200 140098 120000
rect 141606 119200 141662 120000
rect 143170 119200 143226 120000
rect 144734 119200 144790 120000
rect 146298 119200 146354 120000
rect 147862 119200 147918 120000
rect 149426 119200 149482 120000
rect 150990 119200 151046 120000
rect 152554 119200 152610 120000
rect 154118 119200 154174 120000
rect 155682 119200 155738 120000
rect 157246 119200 157302 120000
rect 158810 119200 158866 120000
rect 160374 119200 160430 120000
rect 161938 119200 161994 120000
rect 163502 119200 163558 120000
rect 165066 119200 165122 120000
rect 166630 119200 166686 120000
rect 168194 119200 168250 120000
rect 169758 119200 169814 120000
rect 171322 119200 171378 120000
rect 172886 119200 172942 120000
rect 174450 119200 174506 120000
rect 176014 119200 176070 120000
rect 177578 119200 177634 120000
rect 179142 119200 179198 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148598 0 148654 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168746 0 168802 800
rect 169114 0 169170 800
rect 169482 0 169538 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170586 0 170642 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 112 119144 698 119200
rect 866 119144 2262 119200
rect 2430 119144 3826 119200
rect 3994 119144 5390 119200
rect 5558 119144 6954 119200
rect 7122 119144 8518 119200
rect 8686 119144 10082 119200
rect 10250 119144 11646 119200
rect 11814 119144 13210 119200
rect 13378 119144 14774 119200
rect 14942 119144 16338 119200
rect 16506 119144 17902 119200
rect 18070 119144 19466 119200
rect 19634 119144 21030 119200
rect 21198 119144 22594 119200
rect 22762 119144 24158 119200
rect 24326 119144 25722 119200
rect 25890 119144 27286 119200
rect 27454 119144 28850 119200
rect 29018 119144 30414 119200
rect 30582 119144 31978 119200
rect 32146 119144 33542 119200
rect 33710 119144 35106 119200
rect 35274 119144 36670 119200
rect 36838 119144 38234 119200
rect 38402 119144 39798 119200
rect 39966 119144 41362 119200
rect 41530 119144 42926 119200
rect 43094 119144 44490 119200
rect 44658 119144 46054 119200
rect 46222 119144 47618 119200
rect 47786 119144 49182 119200
rect 49350 119144 50746 119200
rect 50914 119144 52310 119200
rect 52478 119144 53874 119200
rect 54042 119144 55438 119200
rect 55606 119144 57002 119200
rect 57170 119144 58566 119200
rect 58734 119144 60130 119200
rect 60298 119144 61694 119200
rect 61862 119144 63258 119200
rect 63426 119144 64822 119200
rect 64990 119144 66386 119200
rect 66554 119144 67950 119200
rect 68118 119144 69514 119200
rect 69682 119144 71078 119200
rect 71246 119144 72642 119200
rect 72810 119144 74206 119200
rect 74374 119144 75770 119200
rect 75938 119144 77334 119200
rect 77502 119144 78898 119200
rect 79066 119144 80462 119200
rect 80630 119144 82026 119200
rect 82194 119144 83590 119200
rect 83758 119144 85154 119200
rect 85322 119144 86718 119200
rect 86886 119144 88282 119200
rect 88450 119144 89846 119200
rect 90014 119144 91502 119200
rect 91670 119144 93066 119200
rect 93234 119144 94630 119200
rect 94798 119144 96194 119200
rect 96362 119144 97758 119200
rect 97926 119144 99322 119200
rect 99490 119144 100886 119200
rect 101054 119144 102450 119200
rect 102618 119144 104014 119200
rect 104182 119144 105578 119200
rect 105746 119144 107142 119200
rect 107310 119144 108706 119200
rect 108874 119144 110270 119200
rect 110438 119144 111834 119200
rect 112002 119144 113398 119200
rect 113566 119144 114962 119200
rect 115130 119144 116526 119200
rect 116694 119144 118090 119200
rect 118258 119144 119654 119200
rect 119822 119144 121218 119200
rect 121386 119144 122782 119200
rect 122950 119144 124346 119200
rect 124514 119144 125910 119200
rect 126078 119144 127474 119200
rect 127642 119144 129038 119200
rect 129206 119144 130602 119200
rect 130770 119144 132166 119200
rect 132334 119144 133730 119200
rect 133898 119144 135294 119200
rect 135462 119144 136858 119200
rect 137026 119144 138422 119200
rect 138590 119144 139986 119200
rect 140154 119144 141550 119200
rect 141718 119144 143114 119200
rect 143282 119144 144678 119200
rect 144846 119144 146242 119200
rect 146410 119144 147806 119200
rect 147974 119144 149370 119200
rect 149538 119144 150934 119200
rect 151102 119144 152498 119200
rect 152666 119144 154062 119200
rect 154230 119144 155626 119200
rect 155794 119144 157190 119200
rect 157358 119144 158754 119200
rect 158922 119144 160318 119200
rect 160486 119144 161882 119200
rect 162050 119144 163446 119200
rect 163614 119144 165010 119200
rect 165178 119144 166574 119200
rect 166742 119144 168138 119200
rect 168306 119144 169702 119200
rect 169870 119144 171266 119200
rect 171434 119144 172830 119200
rect 172998 119144 174394 119200
rect 174562 119144 175958 119200
rect 176126 119144 177522 119200
rect 177690 119144 179086 119200
rect 179254 119144 179840 119200
rect 112 856 179840 119144
rect 222 800 330 856
rect 498 800 698 856
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4378 856
rect 4546 800 4746 856
rect 4914 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5850 856
rect 6018 800 6218 856
rect 6386 800 6586 856
rect 6754 800 6954 856
rect 7122 800 7322 856
rect 7490 800 7690 856
rect 7858 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8794 856
rect 8962 800 9162 856
rect 9330 800 9530 856
rect 9698 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10634 856
rect 10802 800 11002 856
rect 11170 800 11370 856
rect 11538 800 11738 856
rect 11906 800 12106 856
rect 12274 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13578 856
rect 13746 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15050 856
rect 15218 800 15418 856
rect 15586 800 15786 856
rect 15954 800 16154 856
rect 16322 800 16522 856
rect 16690 800 16890 856
rect 17058 800 17258 856
rect 17426 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18730 856
rect 18898 800 19098 856
rect 19266 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23146 856
rect 23314 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26734 856
rect 26902 800 27102 856
rect 27270 800 27470 856
rect 27638 800 27838 856
rect 28006 800 28206 856
rect 28374 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29310 856
rect 29478 800 29678 856
rect 29846 800 30046 856
rect 30214 800 30414 856
rect 30582 800 30782 856
rect 30950 800 31150 856
rect 31318 800 31518 856
rect 31686 800 31886 856
rect 32054 800 32254 856
rect 32422 800 32622 856
rect 32790 800 32990 856
rect 33158 800 33358 856
rect 33526 800 33726 856
rect 33894 800 34094 856
rect 34262 800 34462 856
rect 34630 800 34830 856
rect 34998 800 35198 856
rect 35366 800 35566 856
rect 35734 800 35934 856
rect 36102 800 36302 856
rect 36470 800 36670 856
rect 36838 800 37038 856
rect 37206 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39614 856
rect 39782 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43294 856
rect 43462 800 43662 856
rect 43830 800 44030 856
rect 44198 800 44398 856
rect 44566 800 44766 856
rect 44934 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45870 856
rect 46038 800 46238 856
rect 46406 800 46606 856
rect 46774 800 46974 856
rect 47142 800 47342 856
rect 47510 800 47710 856
rect 47878 800 48078 856
rect 48246 800 48446 856
rect 48614 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49550 856
rect 49718 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50654 856
rect 50822 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51666 856
rect 51834 800 52034 856
rect 52202 800 52402 856
rect 52570 800 52770 856
rect 52938 800 53138 856
rect 53306 800 53506 856
rect 53674 800 53874 856
rect 54042 800 54242 856
rect 54410 800 54610 856
rect 54778 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55714 856
rect 55882 800 56082 856
rect 56250 800 56450 856
rect 56618 800 56818 856
rect 56986 800 57186 856
rect 57354 800 57554 856
rect 57722 800 57922 856
rect 58090 800 58290 856
rect 58458 800 58658 856
rect 58826 800 59026 856
rect 59194 800 59394 856
rect 59562 800 59762 856
rect 59930 800 60130 856
rect 60298 800 60498 856
rect 60666 800 60866 856
rect 61034 800 61234 856
rect 61402 800 61602 856
rect 61770 800 61970 856
rect 62138 800 62338 856
rect 62506 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63810 856
rect 63978 800 64178 856
rect 64346 800 64546 856
rect 64714 800 64914 856
rect 65082 800 65282 856
rect 65450 800 65650 856
rect 65818 800 66018 856
rect 66186 800 66386 856
rect 66554 800 66754 856
rect 66922 800 67122 856
rect 67290 800 67490 856
rect 67658 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68594 856
rect 68762 800 68962 856
rect 69130 800 69330 856
rect 69498 800 69698 856
rect 69866 800 70066 856
rect 70234 800 70434 856
rect 70602 800 70802 856
rect 70970 800 71170 856
rect 71338 800 71538 856
rect 71706 800 71906 856
rect 72074 800 72274 856
rect 72442 800 72642 856
rect 72810 800 73010 856
rect 73178 800 73378 856
rect 73546 800 73746 856
rect 73914 800 74114 856
rect 74282 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75218 856
rect 75386 800 75586 856
rect 75754 800 75954 856
rect 76122 800 76322 856
rect 76490 800 76690 856
rect 76858 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78806 856
rect 78974 800 79174 856
rect 79342 800 79542 856
rect 79710 800 79910 856
rect 80078 800 80278 856
rect 80446 800 80646 856
rect 80814 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81750 856
rect 81918 800 82118 856
rect 82286 800 82486 856
rect 82654 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83958 856
rect 84126 800 84326 856
rect 84494 800 84694 856
rect 84862 800 85062 856
rect 85230 800 85430 856
rect 85598 800 85798 856
rect 85966 800 86166 856
rect 86334 800 86534 856
rect 86702 800 86902 856
rect 87070 800 87270 856
rect 87438 800 87638 856
rect 87806 800 88006 856
rect 88174 800 88374 856
rect 88542 800 88742 856
rect 88910 800 89110 856
rect 89278 800 89478 856
rect 89646 800 89846 856
rect 90014 800 90214 856
rect 90382 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91686 856
rect 91854 800 92054 856
rect 92222 800 92422 856
rect 92590 800 92790 856
rect 92958 800 93158 856
rect 93326 800 93526 856
rect 93694 800 93894 856
rect 94062 800 94262 856
rect 94430 800 94630 856
rect 94798 800 94998 856
rect 95166 800 95366 856
rect 95534 800 95734 856
rect 95902 800 96102 856
rect 96270 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97206 856
rect 97374 800 97574 856
rect 97742 800 97942 856
rect 98110 800 98310 856
rect 98478 800 98678 856
rect 98846 800 99046 856
rect 99214 800 99414 856
rect 99582 800 99782 856
rect 99950 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101254 856
rect 101422 800 101622 856
rect 101790 800 101990 856
rect 102158 800 102358 856
rect 102526 800 102726 856
rect 102894 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105946 856
rect 106114 800 106314 856
rect 106482 800 106682 856
rect 106850 800 107050 856
rect 107218 800 107418 856
rect 107586 800 107786 856
rect 107954 800 108154 856
rect 108322 800 108522 856
rect 108690 800 108890 856
rect 109058 800 109258 856
rect 109426 800 109626 856
rect 109794 800 109994 856
rect 110162 800 110362 856
rect 110530 800 110730 856
rect 110898 800 111098 856
rect 111266 800 111466 856
rect 111634 800 111834 856
rect 112002 800 112202 856
rect 112370 800 112570 856
rect 112738 800 112938 856
rect 113106 800 113306 856
rect 113474 800 113674 856
rect 113842 800 114042 856
rect 114210 800 114410 856
rect 114578 800 114778 856
rect 114946 800 115146 856
rect 115314 800 115514 856
rect 115682 800 115882 856
rect 116050 800 116250 856
rect 116418 800 116618 856
rect 116786 800 116986 856
rect 117154 800 117354 856
rect 117522 800 117722 856
rect 117890 800 118090 856
rect 118258 800 118458 856
rect 118626 800 118826 856
rect 118994 800 119194 856
rect 119362 800 119562 856
rect 119730 800 119930 856
rect 120098 800 120298 856
rect 120466 800 120666 856
rect 120834 800 121034 856
rect 121202 800 121402 856
rect 121570 800 121770 856
rect 121938 800 122138 856
rect 122306 800 122506 856
rect 122674 800 122874 856
rect 123042 800 123242 856
rect 123410 800 123610 856
rect 123778 800 123978 856
rect 124146 800 124346 856
rect 124514 800 124714 856
rect 124882 800 125082 856
rect 125250 800 125450 856
rect 125618 800 125818 856
rect 125986 800 126186 856
rect 126354 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127290 856
rect 127458 800 127658 856
rect 127826 800 128026 856
rect 128194 800 128394 856
rect 128562 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130510 856
rect 130678 800 130878 856
rect 131046 800 131246 856
rect 131414 800 131614 856
rect 131782 800 131982 856
rect 132150 800 132350 856
rect 132518 800 132718 856
rect 132886 800 133086 856
rect 133254 800 133454 856
rect 133622 800 133822 856
rect 133990 800 134190 856
rect 134358 800 134558 856
rect 134726 800 134926 856
rect 135094 800 135294 856
rect 135462 800 135662 856
rect 135830 800 136030 856
rect 136198 800 136398 856
rect 136566 800 136766 856
rect 136934 800 137134 856
rect 137302 800 137502 856
rect 137670 800 137870 856
rect 138038 800 138238 856
rect 138406 800 138606 856
rect 138774 800 138974 856
rect 139142 800 139342 856
rect 139510 800 139710 856
rect 139878 800 140078 856
rect 140246 800 140446 856
rect 140614 800 140814 856
rect 140982 800 141182 856
rect 141350 800 141550 856
rect 141718 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142654 856
rect 142822 800 143022 856
rect 143190 800 143390 856
rect 143558 800 143758 856
rect 143926 800 144126 856
rect 144294 800 144494 856
rect 144662 800 144862 856
rect 145030 800 145230 856
rect 145398 800 145598 856
rect 145766 800 145966 856
rect 146134 800 146334 856
rect 146502 800 146702 856
rect 146870 800 147070 856
rect 147238 800 147438 856
rect 147606 800 147806 856
rect 147974 800 148174 856
rect 148342 800 148542 856
rect 148710 800 148910 856
rect 149078 800 149278 856
rect 149446 800 149646 856
rect 149814 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150750 856
rect 150918 800 151118 856
rect 151286 800 151486 856
rect 151654 800 151854 856
rect 152022 800 152222 856
rect 152390 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153326 856
rect 153494 800 153694 856
rect 153862 800 154062 856
rect 154230 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160594 856
rect 160762 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162066 856
rect 162234 800 162434 856
rect 162602 800 162802 856
rect 162970 800 163170 856
rect 163338 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164274 856
rect 164442 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166482 856
rect 166650 800 166850 856
rect 167018 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167954 856
rect 168122 800 168322 856
rect 168490 800 168690 856
rect 168858 800 169058 856
rect 169226 800 169426 856
rect 169594 800 169794 856
rect 169962 800 170162 856
rect 170330 800 170530 856
rect 170698 800 170898 856
rect 171066 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173106 856
rect 173274 800 173474 856
rect 173642 800 173842 856
rect 174010 800 174210 856
rect 174378 800 174578 856
rect 174746 800 174946 856
rect 175114 800 175314 856
rect 175482 800 175682 856
rect 175850 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178258 856
rect 178426 800 178626 856
rect 178794 800 178994 856
rect 179162 800 179362 856
rect 179530 800 179730 856
<< metal3 >>
rect 179200 59984 180000 60104
<< obsm3 >>
rect 1669 60184 179200 117537
rect 1669 59904 179120 60184
rect 1669 2143 179200 59904
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 52366 119200 52422 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57058 119200 57114 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 66442 119200 66498 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 71134 119200 71190 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 75826 119200 75882 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 85210 119200 85266 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 94686 119200 94742 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 99378 119200 99434 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 104070 119200 104126 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 113454 119200 113510 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 122838 119200 122894 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 127530 119200 127586 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 132222 119200 132278 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10138 119200 10194 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 141606 119200 141662 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 146298 119200 146354 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 150990 119200 151046 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 165066 119200 165122 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 174450 119200 174506 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14830 119200 14886 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 19522 119200 19578 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 28906 119200 28962 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 33598 119200 33654 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 38290 119200 38346 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 42982 119200 43038 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2318 119200 2374 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 49238 119200 49294 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 63314 119200 63370 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 68006 119200 68062 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 72698 119200 72754 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 77390 119200 77446 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 82082 119200 82138 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 86774 119200 86830 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 91558 119200 91614 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7010 119200 7066 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 100942 119200 100998 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 110326 119200 110382 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 115018 119200 115074 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 124402 119200 124458 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 129094 119200 129150 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 133786 119200 133842 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 138478 119200 138534 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11702 119200 11758 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 143170 119200 143226 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 147862 119200 147918 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 152554 119200 152610 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 157246 119200 157302 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 161938 119200 161994 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 166630 119200 166686 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 171322 119200 171378 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 176014 119200 176070 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 16394 119200 16450 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 21086 119200 21142 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 35162 119200 35218 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 39854 119200 39910 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 50802 119200 50858 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 64878 119200 64934 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 78954 119200 79010 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 83646 119200 83702 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 88338 119200 88394 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 93122 119200 93178 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 119200 8630 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 97814 119200 97870 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 102506 119200 102562 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 116582 119200 116638 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 121274 119200 121330 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 125966 119200 126022 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 130658 119200 130714 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 135350 119200 135406 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 140042 119200 140098 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13266 119200 13322 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 144734 119200 144790 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 149426 119200 149482 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 154118 119200 154174 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 158810 119200 158866 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 163502 119200 163558 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 168194 119200 168250 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 172886 119200 172942 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 17958 119200 18014 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 22650 119200 22706 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 27342 119200 27398 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 32034 119200 32090 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 36726 119200 36782 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 41418 119200 41474 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 46110 119200 46166 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179200 59984 180000 60104 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179142 119200 179198 120000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 169114 0 169170 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 620 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 626 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 627 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 632 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 633 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 638 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 639 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 651 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 652 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 653 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 655 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj.gds
string GDS_END 17323698
string GDS_START 617578
<< end >>

