* NGSPICE file created from user_proj.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

.subckt user_proj io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vccd1 vssd1
+ vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vssa2_uq0 vssa2_uq1 vssa2_uq2 vssa2_uq3 vssa2_uq4
+ vssa1_uq0 vssa1_uq1 vssa1_uq2 vssa1_uq3 vssa1_uq4 vssd2_uq0 vssd2_uq1 vssd2_uq2
+ vssd2_uq3 vssd2_uq4 vdda2_uq0 vdda2_uq1 vdda2_uq2 vdda2_uq3 vdda2_uq4 vdda1_uq0
+ vdda1_uq1 vdda1_uq2 vdda1_uq3 vdda1_uq4 vccd2_uq0 vccd2_uq1 vccd2_uq2 vccd2_uq3
+ vccd2_uq4
XFILLER_136_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2106_ _2185_/A vssd1 vssd1 vccd1 vccd1 _2106_/X sky130_fd_sc_hd__clkbuf_2
X_3086_ _3086_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3086_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ _2037_/A _2053_/B vssd1 vssd1 vccd1 vccd1 _2087_/A sky130_fd_sc_hd__or2_1
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2939_ _3095_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2939_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_178_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1270_ _2199_/A vssd1 vssd1 vccd1 vccd1 _1270_/X sky130_fd_sc_hd__buf_1
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2724_ _2729_/CLK _2724_/D vssd1 vssd1 vccd1 vccd1 _2724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2655_ _1722_/Y _1667_/Y _1807_/Y _1677_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2655_/X sky130_fd_sc_hd__mux4_1
Xoutput401 _2320_/X vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput412 _2745_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput423 _2755_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__clkbuf_2
Xoutput434 _2212_/LO vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__clkbuf_2
X_1606_ _1606_/A _1606_/B vssd1 vssd1 vccd1 vccd1 _1608_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2586_ _2718_/Q _2585_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__mux2_1
Xoutput445 _2216_/LO vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__clkbuf_2
Xoutput456 _2360_/X vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__clkbuf_2
Xoutput467 _2370_/X vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput478 _2230_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__clkbuf_2
X_1537_ _1443_/B _1447_/A _1442_/A _1448_/B vssd1 vssd1 vccd1 vccd1 _1537_/X sky130_fd_sc_hd__o22a_1
Xoutput489 _2240_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1468_ _1468_/A _1468_/B vssd1 vssd1 vccd1 vccd1 _3093_/D sky130_fd_sc_hd__nor2_4
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1399_ _2945_/Q _1371_/X _2984_/Q _1372_/X _1398_/X vssd1 vssd1 vccd1 vccd1 _1399_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3069_ _3108_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3069_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2440_ _2600_/X _2439_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2440_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2371_ _2750_/Q vssd1 vssd1 vccd1 vccd1 _2371_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1322_ _2934_/Q _1303_/X _2973_/Q _1304_/X _1321_/X vssd1 vssd1 vccd1 vccd1 _1322_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_64_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1253_ _3041_/Q _2187_/X _2885_/Q _2188_/X vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2707_ _2722_/CLK _2707_/D vssd1 vssd1 vccd1 vccd1 _2707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2638_ _2191_/X _2803_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2569_ _1994_/X _2726_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1940_ _1940_/A vssd1 vssd1 vccd1 vccd1 _1941_/B sky130_fd_sc_hd__inv_2
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1871_ _1872_/A _2462_/X vssd1 vssd1 vccd1 vccd1 _2704_/D sky130_fd_sc_hd__and2_1
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2423_ _2584_/X _2423_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2354_ _2733_/Q vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__buf_4
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1305_ _3048_/Q _1294_/X _2892_/Q _1295_/X vssd1 vssd1 vccd1 vccd1 _1305_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2285_ vssd1 vssd1 vccd1 vccd1 _2285_/HI _2285_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2088_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2508_/S sky130_fd_sc_hd__or2_1
XFILLER_208_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _3089_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2972_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_206_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1923_ _2671_/Q _1921_/X _2703_/Q _1922_/X vssd1 vssd1 vccd1 vccd1 _2671_/D sky130_fd_sc_hd__a22o_1
XFILLER_148_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1854_ _1854_/A _2426_/X vssd1 vssd1 vccd1 vccd1 _2718_/D sky130_fd_sc_hd__and2_1
XFILLER_15_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1785_ _1783_/X _1784_/X _1783_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2406_ _2566_/X _2405_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2337_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2268_ vssd1 vssd1 vccd1 vccd1 _2268_/HI _2268_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _2199_/A vssd1 vssd1 vccd1 vccd1 _2199_/X sky130_fd_sc_hd__buf_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput301 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input301/X sky130_fd_sc_hd__buf_1
XPHY_7322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput312 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 input312/X sky130_fd_sc_hd__buf_1
XPHY_7333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput323 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 input323/X sky130_fd_sc_hd__buf_1
XPHY_7344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput334 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 _2441_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput345 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 _2429_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput356 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 _2455_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput367 wbs_we_i vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_5 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1570_ _1449_/A _1464_/B _1450_/B _1462_/A vssd1 vssd1 vccd1 vccd1 _1570_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2122_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__inv_2
XFILLER_39_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2053_ _2053_/A _2053_/B vssd1 vssd1 vccd1 vccd1 _2078_/A sky130_fd_sc_hd__or2_1
XFILLER_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2955_ _3111_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2955_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1906_ _2682_/Q _1900_/X _2714_/Q _1901_/X vssd1 vssd1 vccd1 vccd1 _2682_/D sky130_fd_sc_hd__a22o_1
XFILLER_108_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2886_ _3081_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2886_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_178_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1837_ _2650_/X vssd1 vssd1 vccd1 vccd1 _1882_/A sky130_fd_sc_hd__inv_2
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1768_ _1716_/Y _1713_/Y _2795_/Q _2762_/Q vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__a22o_1
XFILLER_89_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1699_ _2780_/Q vssd1 vssd1 vccd1 vccd1 _1699_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput120 la_data_in[58] vssd1 vssd1 vccd1 vccd1 _1483_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput131 la_data_in[68] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__buf_1
XPHY_7152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput142 la_data_in[78] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__buf_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput153 la_data_in[88] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_1
XFILLER_37_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 la_data_in[98] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_1
XPHY_7185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_oenb[107] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__buf_1
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 la_oenb[117] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_hd__buf_1
XPHY_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput197 la_oenb[127] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_1
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2740_ _2761_/CLK _2740_/D vssd1 vssd1 vccd1 vccd1 _2740_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2671_ _2722_/CLK _2671_/D vssd1 vssd1 vccd1 vccd1 _2671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1622_ _1636_/A _1611_/C _2104_/A _1613_/X vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__o31a_4
Xoutput605 _2672_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1553_ _1549_/X _1552_/X _1549_/X _1552_/X vssd1 vssd1 vccd1 vccd1 _1554_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1484_ _1490_/A _1484_/B vssd1 vssd1 vccd1 vccd1 _3100_/D sky130_fd_sc_hd__nor2_4
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2105_ _2105_/A vssd1 vssd1 vccd1 vccd1 _2185_/A sky130_fd_sc_hd__buf_1
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3085_ _3085_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3085_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2036_ _2625_/S _2040_/B vssd1 vssd1 vccd1 vccd1 _2061_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2938_ _3094_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2938_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_143_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2869_ _3103_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2869_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2723_ _2728_/CLK _2723_/D vssd1 vssd1 vccd1 vccd1 _2723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2654_ _2030_/X _2622_/X _2623_/X _2624_/X _2626_/S _2053_/B vssd1 vssd1 vccd1 vccd1
+ _2654_/X sky130_fd_sc_hd__mux4_1
Xoutput402 _2321_/X vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput413 _2746_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1605_ _1605_/A _1605_/B vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__or2_1
Xoutput424 _2756_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__clkbuf_2
Xoutput435 _2213_/LO vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__clkbuf_2
X_2585_ _2006_/X _2718_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__mux2_1
Xoutput446 _2217_/LO vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__clkbuf_2
Xoutput457 _2361_/X vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1536_ _1527_/X _1535_/X _1527_/X _1535_/X vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__o2bb2a_1
Xoutput468 _2371_/X vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__clkbuf_2
Xoutput479 _2231_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1467_ _1467_/A vssd1 vssd1 vccd1 vccd1 _1468_/B sky130_fd_sc_hd__inv_2
XFILLER_25_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1398_ _3062_/Q _1396_/X _2906_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1398_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3068_ _3107_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3068_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _2697_/Q _2557_/S _2018_/Y _2664_/D vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__a22o_1
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2370_ _2749_/Q vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1321_ _3051_/Q _1294_/X _2895_/Q _1295_/X vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__a22o_1
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1252_ _3080_/Q _2185_/X _3002_/Q _2196_/X vssd1 vssd1 vccd1 vccd1 _1252_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2706_ _2722_/CLK _2706_/D vssd1 vssd1 vccd1 vccd1 _2706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2637_ _2183_/X _2802_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2568_ _2725_/Q _2567_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1519_ _1481_/A _1488_/B _1482_/B _1487_/A vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2499_ _2628_/X _2774_/Q _2499_/S vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1870_ _1872_/A _2432_/X vssd1 vssd1 vccd1 vccd1 _2705_/D sky130_fd_sc_hd__and2_1
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2422_ _2582_/X _2421_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2353_ _2732_/Q vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__buf_4
XFILLER_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1304_ _2199_/A vssd1 vssd1 vccd1 vccd1 _1304_/X sky130_fd_sc_hd__buf_1
XFILLER_211_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2284_ vssd1 vssd1 vccd1 vccd1 _2284_/HI _2284_/LO sky130_fd_sc_hd__conb_1
XFILLER_85_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1999_ _2727_/Q _1996_/B _1998_/Y _2728_/Q _1996_/Y vssd1 vssd1 vccd1 vccd1 _1999_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_197_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2971_ _3088_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2971_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_56_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1853_ _1854_/A _2428_/X vssd1 vssd1 vccd1 vccd1 _2719_/D sky130_fd_sc_hd__and2_1
XFILLER_50_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1784_ _2778_/Q _2776_/Q _1714_/Y _1669_/Y vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__o22a_1
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2405_ _2566_/X _2405_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2336_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2267_ vssd1 vssd1 vccd1 vccd1 _2267_/HI _2267_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2198_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2198_/X sky130_fd_sc_hd__buf_1
XFILLER_26_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput302 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input302/X sky130_fd_sc_hd__buf_1
XPHY_7323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput313 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 input313/X sky130_fd_sc_hd__buf_1
XFILLER_0_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput324 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 input324/X sky130_fd_sc_hd__buf_1
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput335 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 _2443_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput346 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 _2399_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput357 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 _2457_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_6 _1398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2121_ _2121_/A _2397_/S _2396_/S vssd1 vssd1 vccd1 vccd1 _2122_/A sky130_fd_sc_hd__or3_4
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2052_ _2060_/A _2077_/A vssd1 vssd1 vccd1 vccd1 _2481_/S sky130_fd_sc_hd__or2_1
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2954_ _3110_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2954_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1905_ _2683_/Q _1900_/X _2715_/Q _1901_/X vssd1 vssd1 vccd1 vccd1 _2683_/D sky130_fd_sc_hd__a22o_1
XFILLER_143_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2885_ _3080_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2885_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1836_ _1742_/B _1836_/B _1932_/B vssd1 vssd1 vccd1 vccd1 _2729_/D sky130_fd_sc_hd__and3b_2
XFILLER_102_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1767_ _2790_/Q _2793_/Q _1705_/Y _2030_/A vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__o22a_1
XFILLER_89_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1698_ _2764_/Q vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2319_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 la_data_in[49] vssd1 vssd1 vccd1 vccd1 _1462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput121 la_data_in[59] vssd1 vssd1 vccd1 vccd1 _1485_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput132 la_data_in[69] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__buf_1
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput143 la_data_in[79] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__buf_1
XPHY_7164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 la_data_in[89] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__buf_1
XPHY_7175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput165 la_data_in[99] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_1
XPHY_7186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 la_oenb[108] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_hd__buf_1
XPHY_7197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput187 la_oenb[118] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_hd__buf_1
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput198 la_oenb[12] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__buf_1
XFILLER_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2670_ _2722_/CLK _2670_/D vssd1 vssd1 vccd1 vccd1 _2670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1621_ _1636_/A _1617_/B _2398_/X _1618_/X _1879_/A vssd1 vssd1 vccd1 vccd1 _1621_/X
+ sky130_fd_sc_hd__o41a_4
Xoutput606 _2673_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1552_ _1437_/B _1551_/A _1436_/A _1551_/Y vssd1 vssd1 vccd1 vccd1 _1552_/X sky130_fd_sc_hd__o22a_1
XFILLER_181_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1483_ _1483_/A vssd1 vssd1 vccd1 vccd1 _1484_/B sky130_fd_sc_hd__inv_2
XFILLER_141_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2104_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__inv_2
XFILLER_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3084_ _3084_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3084_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2035_ _2047_/A _2086_/A vssd1 vssd1 vccd1 vccd1 _2463_/S sky130_fd_sc_hd__or2_1
XFILLER_130_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2937_ _3093_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2937_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2868_ _3102_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2868_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1819_ _1731_/Y _1765_/X _1731_/Y _1765_/X vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2799_ _2799_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2799_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_163_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2722_ _2722_/CLK _2722_/D vssd1 vssd1 vccd1 vccd1 _2722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653_ _2653_/A0 _2653_/A1 _2653_/S vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__mux2_8
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput403 _2322_/X vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_145_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput414 _2747_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__clkbuf_2
X_1604_ _1605_/A _1605_/B vssd1 vssd1 vccd1 vccd1 _1606_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput425 _2757_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__clkbuf_2
X_2584_ _2717_/Q _2583_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput436 _2214_/LO vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__clkbuf_2
Xoutput447 _2218_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput458 _2228_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__clkbuf_2
X_1535_ _1492_/B _1534_/X _1492_/B _1534_/X vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__a2bb2o_1
Xoutput469 _2229_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1466_ _1468_/A _1466_/B vssd1 vssd1 vccd1 vccd1 _3092_/D sky130_fd_sc_hd__nor2_4
XFILLER_29_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1397_ _2123_/A vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__buf_1
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3067_ _3106_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3067_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_58_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2018_ _2697_/Q vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1320_ _3090_/Q _1292_/X _3012_/Q _1301_/X vssd1 vssd1 vccd1 vccd1 _1320_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1251_ _2134_/A _2641_/X _1494_/A vssd1 vssd1 vccd1 vccd1 _2767_/D sky130_fd_sc_hd__a21o_1
XFILLER_133_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2705_ _2722_/CLK _2705_/D vssd1 vssd1 vccd1 vccd1 _2705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2636_ _2177_/X _2801_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2567_ _1991_/X _2725_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1518_ _1470_/A _1486_/B _1471_/B _1485_/A vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2498_ _2497_/X _2773_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1449_ _1449_/A vssd1 vssd1 vccd1 vccd1 _1450_/B sky130_fd_sc_hd__inv_2
XFILLER_64_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2421_ _2582_/X _2421_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2421_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2352_ _2731_/Q vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__buf_4
XFILLER_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1303_ _2198_/A vssd1 vssd1 vccd1 vccd1 _1303_/X sky130_fd_sc_hd__buf_1
X_2283_ vssd1 vssd1 vccd1 vccd1 _2283_/HI _2283_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1998_ _2728_/Q vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2619_ _2703_/Q _2618_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2970_ _3087_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2970_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1921_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1852_ _1854_/A _2430_/X vssd1 vssd1 vccd1 vccd1 _2720_/D sky130_fd_sc_hd__and2_1
XFILLER_54_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1783_ _1709_/Y _1782_/X _1709_/Y _1782_/X vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2404_ _2564_/X _2403_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2404_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2335_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2266_ vssd1 vssd1 vccd1 vccd1 _2266_/HI _2266_/LO sky130_fd_sc_hd__conb_1
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2197_ _3077_/Q _2185_/X _2999_/Q _2196_/X vssd1 vssd1 vccd1 vccd1 _2197_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput303 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input303/X sky130_fd_sc_hd__buf_1
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput314 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 input314/X sky130_fd_sc_hd__buf_1
XPHY_7335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput325 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 input325/X sky130_fd_sc_hd__buf_1
XPHY_7346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput336 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 _2445_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput347 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 _2401_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput358 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 _2459_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 _2664_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2120_ _2187_/A vssd1 vssd1 vccd1 vccd1 _2120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2051_ _2059_/A _2073_/A vssd1 vssd1 vccd1 vccd1 _2077_/A sky130_fd_sc_hd__or2_1
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2953_ _3109_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2953_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1904_ _2684_/Q _1900_/X _2716_/Q _1901_/X vssd1 vssd1 vccd1 vccd1 _2684_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2884_ _3079_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2884_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_206_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1835_ _2087_/C _2054_/B _2065_/A vssd1 vssd1 vccd1 vccd1 _1932_/B sky130_fd_sc_hd__or3_4
XFILLER_204_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1766_ _1723_/X _1765_/X _1723_/X _1765_/X vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1697_ _2793_/Q vssd1 vssd1 vccd1 vccd1 _2030_/A sky130_fd_sc_hd__inv_2
XFILLER_172_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2318_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2318_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2249_ vssd1 vssd1 vccd1 vccd1 _2249_/HI _2249_/LO sky130_fd_sc_hd__conb_1
XFILLER_187_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _2398_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput111 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _2396_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput122 la_data_in[5] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__buf_1
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 la_data_in[6] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__buf_1
Xinput144 la_data_in[7] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__buf_1
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_data_in[8] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__buf_1
XPHY_7176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_data_in[9] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_1
XPHY_7187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 la_oenb[109] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__buf_1
XFILLER_40_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput188 la_oenb[119] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__buf_1
XPHY_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 la_oenb[13] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__buf_1
XFILLER_40_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1620_ _1636_/A _1617_/B _2397_/X _1618_/X _1879_/A vssd1 vssd1 vccd1 vccd1 _1620_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_138_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput607 _2674_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1551_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1551_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1482_ _1490_/A _1482_/B vssd1 vssd1 vccd1 vccd1 _3099_/D sky130_fd_sc_hd__nor2_4
XFILLER_64_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2103_ _2107_/A _2111_/B vssd1 vssd1 vccd1 vccd1 _2104_/A sky130_fd_sc_hd__or2_2
XFILLER_95_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3083_ _3083_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3083_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2034_ _2065_/A _2059_/A vssd1 vssd1 vccd1 vccd1 _2086_/A sky130_fd_sc_hd__or2_1
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2936_ _3092_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2936_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2867_ _3101_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2867_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1818_ _1818_/A vssd1 vssd1 vccd1 vccd1 _1834_/A sky130_fd_sc_hd__buf_1
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2798_ _2798_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2798_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1749_ _1735_/X _1748_/X _1735_/X _1748_/X vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2721_ _2722_/CLK _2721_/D vssd1 vssd1 vccd1 vccd1 _2721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _1318_/X _2816_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1603_ _1508_/X _1602_/X _1508_/X _1602_/X vssd1 vssd1 vccd1 vccd1 _1605_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput404 _2323_/X vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput415 _2748_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2583_ _2005_/X _2717_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__mux2_1
Xoutput426 _2758_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput437 _2733_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput448 _2352_/X vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1534_ _1427_/B _1428_/A _1426_/A _1429_/B vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput459 _2362_/X vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1465_ _1465_/A vssd1 vssd1 vccd1 vccd1 _1466_/B sky130_fd_sc_hd__inv_2
XFILLER_29_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1396_ _2119_/A vssd1 vssd1 vccd1 vccd1 _1396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3066_ _3105_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3066_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2017_ _2712_/Q _1959_/B _1960_/A vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2919_ _3075_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2919_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1250_ _2650_/X vssd1 vssd1 vccd1 vccd1 _1494_/A sky130_fd_sc_hd__buf_4
XFILLER_172_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2704_ _2722_/CLK _2704_/D vssd1 vssd1 vccd1 vccd1 _2704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2635_ _2172_/X _2839_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2566_ _2724_/Q _2565_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1517_ _1425_/B _1429_/B _1424_/A _1428_/A vssd1 vssd1 vccd1 vccd1 _1517_/X sky130_fd_sc_hd__a22o_1
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2497_ _2496_/X _2773_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1448_ _1456_/A _1448_/B vssd1 vssd1 vccd1 vccd1 _3084_/D sky130_fd_sc_hd__nor2_4
XFILLER_116_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1379_ _3059_/Q _1362_/X _2903_/Q _1363_/X vssd1 vssd1 vccd1 vccd1 _1379_/X sky130_fd_sc_hd__a22o_1
XFILLER_151_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3049_ _3088_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3049_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2420_ _2580_/X _2419_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2351_ _2730_/Q vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__buf_4
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1302_ _3087_/Q _1292_/X _3009_/Q _1301_/X vssd1 vssd1 vccd1 vccd1 _1302_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2282_ vssd1 vssd1 vccd1 vccd1 _2282_/HI _2282_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2727_/Q _1996_/B _1996_/Y vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2618_ _2027_/X _2703_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2549_ _2548_/X _2790_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1920_ _2672_/Q _1914_/X _2704_/Q _1915_/X vssd1 vssd1 vccd1 vccd1 _2672_/D sky130_fd_sc_hd__a22o_1
XFILLER_182_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1851_ _1854_/A _2400_/X vssd1 vssd1 vccd1 vccd1 _2721_/D sky130_fd_sc_hd__and2_1
XFILLER_175_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1782_ _1728_/Y _2781_/Q _2785_/Q _1733_/Y vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__o22a_1
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2403_ _2564_/X _2403_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2403_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2334_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2265_ vssd1 vssd1 vccd1 vccd1 _2265_/HI _2265_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2196_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2196_/X sky130_fd_sc_hd__buf_1
XFILLER_211_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput304 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 input304/X sky130_fd_sc_hd__buf_1
XPHY_7325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput315 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 input315/X sky130_fd_sc_hd__buf_1
XFILLER_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput326 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 input326/X sky130_fd_sc_hd__buf_1
XFILLER_44_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput337 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 _2415_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput348 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 _2403_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput359 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 _2461_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_8 _2944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2050_ _2060_/A _2076_/A vssd1 vssd1 vccd1 vccd1 _2478_/S sky130_fd_sc_hd__or2_1
XFILLER_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _3108_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2952_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1903_ _2685_/Q _1900_/X _2717_/Q _1901_/X vssd1 vssd1 vccd1 vccd1 _2685_/D sky130_fd_sc_hd__a22o_1
XFILLER_203_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2883_ _3078_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2883_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1834_ _1834_/A _2053_/B vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1765_ _2778_/Q _1676_/Y _1714_/Y _2786_/Q vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1696_ _1694_/Y _2799_/Q _2774_/Q _1695_/Y vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__o22a_1
XFILLER_176_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2317_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ vssd1 vssd1 vccd1 vccd1 _2248_/HI _2248_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2179_ _2203_/A _2184_/B _2636_/X vssd1 vssd1 vccd1 vccd1 _2762_/D sky130_fd_sc_hd__and3_1
XFILLER_96_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput101 la_data_in[40] vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__buf_1
XFILLER_81_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput112 la_data_in[50] vssd1 vssd1 vccd1 vccd1 _1465_/A sky130_fd_sc_hd__buf_1
XPHY_7133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 la_data_in[60] vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput134 la_data_in[70] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__buf_1
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 la_data_in[80] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__buf_1
XPHY_7166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 la_data_in[90] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__buf_1
XFILLER_44_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput167 la_oenb[0] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__buf_1
XPHY_7188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput178 la_oenb[10] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__buf_1
XPHY_7199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_oenb[11] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_hd__buf_1
XFILLER_40_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1550_ _1468_/B _1476_/A _1467_/A _1477_/B vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__o22a_1
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1481_ _1481_/A vssd1 vssd1 vccd1 vccd1 _1482_/B sky130_fd_sc_hd__inv_2
XFILLER_113_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2102_ _2102_/A vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__buf_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3082_ _3082_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3082_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_23_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2033_ _2033_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__or2_1
XFILLER_3_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2935_ _3091_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2935_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2866_ _3100_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2866_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1817_ _1832_/A _2053_/A vssd1 vssd1 vccd1 vccd1 _1818_/A sky130_fd_sc_hd__or2_1
X_2797_ _2797_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2797_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1748_ _1673_/Y _1684_/Y _2765_/Q _2763_/Q vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1679_ _1677_/Y _2766_/Q _2770_/Q _1678_/Y vssd1 vssd1 vccd1 vccd1 _1679_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ _2722_/CLK _2720_/D vssd1 vssd1 vccd1 vccd1 _2720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2651_ _1313_/X _2815_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1602_ _1473_/B _1601_/Y _1473_/B _1601_/Y vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput405 _2324_/X vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2582_ _2716_/Q _2581_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput416 _2749_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput427 _2759_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput438 _2734_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__clkbuf_2
X_1533_ _1582_/A _1533_/B vssd1 vssd1 vccd1 vccd1 _3107_/D sky130_fd_sc_hd__nor2_4
XFILLER_86_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput449 _2353_/X vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1464_ _1468_/A _1464_/B vssd1 vssd1 vccd1 vccd1 _3091_/D sky130_fd_sc_hd__nor2_4
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1395_ _3101_/Q _1394_/X _3023_/Q _1369_/X vssd1 vssd1 vccd1 vccd1 _1395_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3065_ _3104_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3065_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2016_ _2711_/Q _1957_/B _1958_/A vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2918_ _3074_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2918_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2849_ _3083_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2849_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2703_ _2722_/CLK _2703_/D vssd1 vssd1 vccd1 vccd1 _2703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2634_ _2167_/X _2838_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2565_ _1988_/X _2724_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1516_ _1516_/A _1582_/A vssd1 vssd1 vccd1 vccd1 _3106_/D sky130_fd_sc_hd__nor2_4
XFILLER_138_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2496_ _2628_/X _2773_/Q _2496_/S vssd1 vssd1 vccd1 vccd1 _2496_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1447_ _1447_/A vssd1 vssd1 vccd1 vccd1 _1448_/B sky130_fd_sc_hd__inv_2
XFILLER_155_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1378_ _3098_/Q _1360_/X _3020_/Q _1369_/X vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3048_ _3087_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3048_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_97_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2350_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1301_ _2196_/A vssd1 vssd1 vccd1 vccd1 _1301_/X sky130_fd_sc_hd__buf_1
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2281_ vssd1 vssd1 vccd1 vccd1 _2281_/HI _2281_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1996_ _2727_/Q _1996_/B vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2617_ _2702_/Q _2616_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2548_ _2547_/X _2790_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ _2478_/X _2767_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__mux2_1
XPHY_6806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1850_ _1854_/A _2402_/X vssd1 vssd1 vccd1 vccd1 _2722_/D sky130_fd_sc_hd__and2_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1781_ _1779_/X _1780_/X _1779_/X _1780_/X vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2402_ _2562_/X _2401_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2402_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2333_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2264_ vssd1 vssd1 vccd1 vccd1 _2264_/HI _2264_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2195_ _2195_/A vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__buf_1
XFILLER_187_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1979_ _1979_/A _2020_/A vssd1 vssd1 vccd1 vccd1 _2413_/S sky130_fd_sc_hd__and2_4
XFILLER_120_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput305 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 input305/X sky130_fd_sc_hd__buf_1
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput316 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 input316/X sky130_fd_sc_hd__buf_1
XPHY_7337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput327 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 input327/X sky130_fd_sc_hd__buf_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput338 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 _2417_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput349 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 _2405_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_9 _2945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2951_ _3107_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2951_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1902_ _2686_/Q _1900_/X _2718_/Q _1901_/X vssd1 vssd1 vccd1 vccd1 _2686_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2882_ _3077_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2882_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1833_ _1833_/A vssd1 vssd1 vccd1 vccd1 _2053_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1764_ _1762_/X _1763_/X _1762_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1695_ _2799_/Q vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2316_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2316_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ vssd1 vssd1 vccd1 vccd1 _2247_/HI _2247_/LO sky130_fd_sc_hd__conb_1
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2178_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2203_/A sky130_fd_sc_hd__buf_1
XFILLER_187_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput102 la_data_in[41] vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__buf_1
XFILLER_27_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 la_data_in[51] vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput124 la_data_in[61] vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput135 la_data_in[71] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__buf_1
XPHY_7156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 la_data_in[81] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__buf_1
XFILLER_44_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_data_in[91] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__buf_1
XPHY_7178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_oenb[100] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__buf_1
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput179 la_oenb[110] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__buf_1
XPHY_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1480_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__buf_4
XFILLER_190_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2101_ _2156_/A vssd1 vssd1 vccd1 vccd1 _2102_/A sky130_fd_sc_hd__buf_1
XFILLER_23_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3081_ _3081_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3081_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2032_ _2054_/B vssd1 vssd1 vccd1 vccd1 _2047_/A sky130_fd_sc_hd__buf_1
XFILLER_97_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2934_ _3090_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2934_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2865_ _3099_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2865_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1816_ _2037_/A vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__inv_2
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2796_ _2796_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2796_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_117_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1747_ _2790_/Q _1713_/Y _1705_/Y _2762_/Q vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1678_ _2766_/Q vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2650_ _2650_/A0 _2650_/A1 _2650_/S vssd1 vssd1 vccd1 vccd1 _2650_/X sky130_fd_sc_hd__mux2_8
XFILLER_200_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1601_ _1591_/X _1600_/X _1591_/X _1600_/X vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_103_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2581_ _2004_/X _2716_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__mux2_1
Xoutput406 _2730_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput417 _2731_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput428 _2732_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput439 _2735_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1532_ _1525_/Y _1531_/Y _1525_/Y _1531_/Y vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_138_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1463_ _1463_/A vssd1 vssd1 vccd1 vccd1 _1464_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1394_ _2105_/A vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__buf_1
XFILLER_132_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3064_ _3103_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3064_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_97_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2015_ _2710_/Q _1955_/B _1956_/A vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _3112_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2917_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_71_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2848_ _3082_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2848_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2779_ _2779_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2779_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_12_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2702_ _2722_/CLK _2702_/D vssd1 vssd1 vccd1 vccd1 _2702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2633_ _2153_/X _2837_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2564_ _2723_/Q _2563_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1515_ _2650_/X _1617_/B vssd1 vssd1 vccd1 vccd1 _1582_/A sky130_fd_sc_hd__or2_4
XFILLER_173_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2495_ _2494_/X _2772_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2495_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1446_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1456_/A sky130_fd_sc_hd__buf_4
XFILLER_190_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1377_ _1387_/A _1401_/B _2387_/X vssd1 vssd1 vccd1 vccd1 _2785_/D sky130_fd_sc_hd__and3_1
XFILLER_56_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3047_ _3086_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3047_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_208_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1300_ _2195_/A vssd1 vssd1 vccd1 vccd1 _1300_/X sky130_fd_sc_hd__buf_1
XFILLER_65_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2280_ vssd1 vssd1 vccd1 vccd1 _2280_/HI _2280_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1995_ _1995_/A vssd1 vssd1 vccd1 vccd1 _1996_/B sky130_fd_sc_hd__inv_2
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2616_ _2026_/X _2702_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2547_ _2628_/X _2790_/Q _2547_/S vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2478_ _2628_/X _2767_/Q _2478_/S vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ _1433_/A _1429_/B vssd1 vssd1 vccd1 vccd1 _3076_/D sky130_fd_sc_hd__nor2_4
XPHY_6829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ _1694_/Y _2783_/Q _2774_/Q _1725_/Y vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__o22a_1
XFILLER_204_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2401_ _2562_/X _2401_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2401_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2332_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2263_ vssd1 vssd1 vccd1 vccd1 _2263_/HI _2263_/LO sky130_fd_sc_hd__conb_1
XFILLER_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2194_ _2203_/A _2203_/B _2638_/X vssd1 vssd1 vccd1 vccd1 _2764_/D sky130_fd_sc_hd__and3_1
XFILLER_61_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1978_ _2721_/Q _1977_/B _1980_/A vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput306 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 input306/X sky130_fd_sc_hd__buf_1
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput317 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input317/X sky130_fd_sc_hd__buf_1
XFILLER_44_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput328 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 input328/X sky130_fd_sc_hd__buf_1
XFILLER_9_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput339 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 _2419_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2950_ _3106_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2950_/Q sky130_fd_sc_hd__dlxtn_1
X_1901_ _1901_/A vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__buf_1
XFILLER_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2881_ _3076_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2881_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ _1832_/A _1832_/B vssd1 vssd1 vccd1 vccd1 _1833_/A sky130_fd_sc_hd__or2_1
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1763_ _2764_/Q _2765_/Q _1698_/Y _1673_/Y vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1694_ _2774_/Q vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2315_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__buf_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2246_ vssd1 vssd1 vccd1 vccd1 _2246_/HI _2246_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2177_ _2840_/Q _2157_/X _2174_/X _2176_/X vssd1 vssd1 vccd1 vccd1 _2177_/X sky130_fd_sc_hd__a211o_1
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput103 la_data_in[42] vssd1 vssd1 vccd1 vccd1 _1447_/A sky130_fd_sc_hd__buf_1
XFILLER_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput114 la_data_in[52] vssd1 vssd1 vccd1 vccd1 _1470_/A sky130_fd_sc_hd__buf_1
XPHY_7135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 la_data_in[62] vssd1 vssd1 vccd1 vccd1 _1491_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 la_data_in[72] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__buf_1
XPHY_7157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput147 la_data_in[82] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__buf_1
XPHY_7168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_data_in[92] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__buf_1
XPHY_7179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput169 la_oenb[101] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__buf_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2100_ _2100_/A vssd1 vssd1 vccd1 vccd1 _2156_/A sky130_fd_sc_hd__inv_2
XFILLER_114_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3080_ _3080_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3080_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_62_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2031_ _2654_/X _2627_/S _1834_/A vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__or3b_1
XFILLER_208_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2933_ _3089_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2933_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2864_ _3098_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2864_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1815_ _1805_/Y _1814_/Y _1805_/Y _1814_/Y vssd1 vssd1 vccd1 vccd1 _2037_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2795_ _2795_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2795_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_30_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1746_ _1746_/A vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__buf_1
XFILLER_85_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1677_ _2770_/Q vssd1 vssd1 vccd1 vccd1 _1677_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ vssd1 vssd1 vccd1 vccd1 _2229_/HI _2229_/LO sky130_fd_sc_hd__conb_1
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1600_ _1592_/X _1599_/Y _1592_/X _1599_/Y vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2580_ _2715_/Q _2579_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput407 _2740_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput418 _2750_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1531_ _1526_/X _1530_/X _1526_/X _1530_/X vssd1 vssd1 vccd1 vccd1 _1531_/Y sky130_fd_sc_hd__a2bb2oi_1
Xoutput429 _2760_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1462_ _1462_/A vssd1 vssd1 vccd1 vccd1 _1463_/A sky130_fd_sc_hd__inv_2
XFILLER_190_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1393_ _1417_/A _1401_/B _2390_/X vssd1 vssd1 vccd1 vccd1 _2788_/D sky130_fd_sc_hd__and3_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3063_ _3102_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3063_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_114_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2014_ _2709_/Q _1953_/B _1954_/A vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2916_ _3111_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2916_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2847_ _3081_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2847_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2778_ _2778_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2778_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_30_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1729_ _2777_/Q _2785_/Q _1727_/Y _1728_/Y vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__o22a_1
XFILLER_156_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2701_ _2722_/CLK _2701_/D vssd1 vssd1 vccd1 vccd1 _2701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2632_ _2145_/X _2836_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2563_ _1985_/X _2723_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1514_ _1609_/B vssd1 vssd1 vccd1 vccd1 _1617_/B sky130_fd_sc_hd__inv_2
X_2494_ _2493_/X _2772_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1445_ _1445_/A _1445_/B vssd1 vssd1 vccd1 vccd1 _3083_/D sky130_fd_sc_hd__nor2_4
XFILLER_136_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1376_ _2193_/A vssd1 vssd1 vccd1 vccd1 _1401_/B sky130_fd_sc_hd__buf_1
XFILLER_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3046_ _3085_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3046_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1994_ _2726_/Q _1993_/B _1995_/A vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2615_ _2701_/Q _2614_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2546_ _2545_/X _2789_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2477_ _2476_/X _2766_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ _1428_/A vssd1 vssd1 vccd1 vccd1 _1429_/B sky130_fd_sc_hd__inv_2
XFILLER_9_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1359_ _1387_/A _1367_/B _2385_/X vssd1 vssd1 vccd1 vccd1 _2783_/D sky130_fd_sc_hd__and3_1
XFILLER_205_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _3107_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3029_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput590 _2687_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2400_ _2560_/X _2399_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2400_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2331_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2262_ vssd1 vssd1 vccd1 vccd1 _2262_/HI _2262_/LO sky130_fd_sc_hd__conb_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2193_ _2193_/A vssd1 vssd1 vccd1 vccd1 _2203_/B sky130_fd_sc_hd__buf_1
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1977_ _2721_/Q _1977_/B vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2529_ _2628_/X _2784_/Q _2529_/S vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput307 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 input307/X sky130_fd_sc_hd__buf_1
XFILLER_48_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput318 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input318/X sky130_fd_sc_hd__buf_1
XPHY_7339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput329 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _1880_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1900_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1900_/X sky130_fd_sc_hd__buf_1
X_2880_ _3075_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2880_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _1821_/Y _1830_/X _1821_/Y _1830_/X vssd1 vssd1 vccd1 vccd1 _1832_/B sky130_fd_sc_hd__o2bb2a_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1762_ _1754_/X _1761_/X _1754_/X _1761_/X vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1693_ _1689_/Y _1692_/X _1689_/Y _1692_/X vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2314_ vssd1 vssd1 vccd1 vccd1 _2314_/HI _2314_/LO sky130_fd_sc_hd__conb_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2245_ vssd1 vssd1 vccd1 vccd1 _2245_/HI _2245_/LO sky130_fd_sc_hd__conb_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2176_ _2918_/Q _2162_/X _2957_/Q _2164_/X _2175_/X vssd1 vssd1 vccd1 vccd1 _2176_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput104 la_data_in[43] vssd1 vssd1 vccd1 vccd1 _1449_/A sky130_fd_sc_hd__buf_1
XPHY_7125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput115 la_data_in[53] vssd1 vssd1 vccd1 vccd1 _1472_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput126 la_data_in[63] vssd1 vssd1 vccd1 vccd1 _1493_/A sky130_fd_sc_hd__buf_2
XPHY_7147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput137 la_data_in[73] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__buf_1
XPHY_7158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 la_data_in[83] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_1
XPHY_7169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput159 la_data_in[93] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__buf_1
XPHY_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2030_ _2030_/A _2625_/S vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__or2_1
XFILLER_149_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2932_ _3088_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2932_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2863_ _3097_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2863_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1814_ _1809_/X _1813_/Y _1809_/X _1813_/Y vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_30_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2794_ _2794_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2794_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1745_ _1832_/A vssd1 vssd1 vccd1 vccd1 _2045_/A sky130_fd_sc_hd__buf_2
XFILLER_201_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1676_ _2786_/Q vssd1 vssd1 vccd1 vccd1 _1676_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ vssd1 vssd1 vccd1 vccd1 _2228_/HI _2228_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _2196_/A vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__buf_1
XFILLER_76_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput408 _2741_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput419 _2751_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1530_ _1528_/X _1529_/X _1528_/X _1529_/X vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1461_ _1468_/A _1461_/B vssd1 vssd1 vccd1 vccd1 _3090_/D sky130_fd_sc_hd__nor2_4
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1392_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__buf_1
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3062_ _3101_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3062_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2013_ _2708_/Q _1951_/B _1952_/A vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__o21a_1
XFILLER_209_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2915_ _3110_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2915_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_56_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2846_ _3080_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2846_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_121_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2777_ _2777_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2777_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1728_ _2785_/Q vssd1 vssd1 vccd1 vccd1 _1728_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1659_ _1659_/A _2480_/X vssd1 vssd1 vccd1 vccd1 _2735_/D sky130_fd_sc_hd__and2_1
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2700_ _2722_/CLK _2700_/D vssd1 vssd1 vccd1 vccd1 _2700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2631_ _2138_/X _2835_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2562_ _2722_/Q _2561_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2562_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1513_ _1500_/X _1512_/X _1500_/X _1512_/X vssd1 vssd1 vccd1 vccd1 _1516_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2493_ _2628_/X _2772_/Q _2493_/S vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1444_ _1527_/A vssd1 vssd1 vccd1 vccd1 _1445_/B sky130_fd_sc_hd__inv_2
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1375_ _2863_/Q _1368_/X _1370_/X _1374_/X vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__a211o_1
XFILLER_136_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3045_ _3084_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3045_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2829_ _3102_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2829_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1993_ _2726_/Q _1993_/B vssd1 vssd1 vccd1 vccd1 _1995_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2614_ _2025_/X _2701_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2545_ _2544_/X _2789_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2476_ _2475_/X _2766_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1427_ _1433_/A _1427_/B vssd1 vssd1 vccd1 vccd1 _3075_/D sky130_fd_sc_hd__nor2_4
XFILLER_25_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1358_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1387_/A sky130_fd_sc_hd__buf_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1289_ _2851_/Q _1266_/X _1286_/X _1288_/X vssd1 vssd1 vccd1 vccd1 _1289_/X sky130_fd_sc_hd__a211o_1
XFILLER_77_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3028_ _3106_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3028_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput580 _2678_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput591 _2688_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2330_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2261_ vssd1 vssd1 vccd1 vccd1 _2261_/HI _2261_/LO sky130_fd_sc_hd__conb_1
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2192_ _2192_/A vssd1 vssd1 vccd1 vccd1 _2193_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1976_ _1976_/A vssd1 vssd1 vccd1 vccd1 _1977_/B sky130_fd_sc_hd__inv_2
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2528_ _2527_/X _2783_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2528_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput308 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 input308/X sky130_fd_sc_hd__buf_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2459_ _2619_/X _2459_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__mux2_1
Xinput319 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 input319/X sky130_fd_sc_hd__buf_1
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _1826_/X _1829_/X _1826_/X _1829_/X vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ _1694_/Y _2782_/Q _2774_/Q _1706_/Y vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__o22a_1
XFILLER_129_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1692_ _2792_/Q _2788_/Q _1746_/A _1691_/Y vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2313_ vssd1 vssd1 vccd1 vccd1 _2313_/HI _2313_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2244_ vssd1 vssd1 vccd1 vccd1 _2244_/HI _2244_/LO sky130_fd_sc_hd__conb_1
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2175_ _3035_/Q _2149_/X _2879_/Q _2150_/X vssd1 vssd1 vccd1 vccd1 _2175_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1959_ _2712_/Q _1959_/B vssd1 vssd1 vccd1 vccd1 _1960_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput105 la_data_in[44] vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__buf_1
XPHY_7126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput116 la_data_in[54] vssd1 vssd1 vccd1 vccd1 _1474_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 la_data_in[64] vssd1 vssd1 vccd1 vccd1 _2653_/A0 sky130_fd_sc_hd__clkbuf_2
XPHY_7148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput138 la_data_in[74] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__buf_1
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 la_data_in[84] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__buf_1
XPHY_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2931_ _3087_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2931_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2862_ _3096_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2862_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1813_ _1810_/X _1812_/Y _1810_/X _1812_/Y vssd1 vssd1 vccd1 vccd1 _1813_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_125_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2793_ _2793_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2793_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_89_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1744_ _2607_/S vssd1 vssd1 vccd1 vccd1 _1832_/A sky130_fd_sc_hd__inv_2
XFILLER_195_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1675_ _2798_/Q _2800_/Q _2798_/Q _2800_/Q vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_85_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2227_ vssd1 vssd1 vccd1 vccd1 _2227_/HI _2227_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2158_ _2158_/A vssd1 vssd1 vccd1 vccd1 _2196_/A sky130_fd_sc_hd__buf_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2089_ _2089_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2556_/S sky130_fd_sc_hd__or2_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput409 _2742_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1460_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1461_/B sky130_fd_sc_hd__inv_2
XFILLER_9_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1391_ _2866_/Q _1368_/X _1388_/X _1390_/X vssd1 vssd1 vccd1 vccd1 _1391_/X sky130_fd_sc_hd__a211o_1
XFILLER_136_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3061_ _3100_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3061_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_7490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2012_ _2707_/Q _1949_/B _1950_/A vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2914_ _3109_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2914_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_56_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2845_ _3079_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2845_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2776_ _2776_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2776_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_89_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1727_ _2777_/Q vssd1 vssd1 vccd1 vccd1 _1727_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1658_ _1659_/A _2483_/X vssd1 vssd1 vccd1 vccd1 _2736_/D sky130_fd_sc_hd__and2_1
XFILLER_67_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1589_ _1440_/A _1527_/X _1441_/B _1445_/B vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__o22a_1
XFILLER_119_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2630_ _2133_/X _2834_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2630_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2561_ _1982_/X _2722_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1512_ _1505_/X _1511_/X _1505_/X _1511_/X vssd1 vssd1 vccd1 vccd1 _1512_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2492_ _2491_/X _2771_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1443_ _1445_/A _1443_/B vssd1 vssd1 vccd1 vccd1 _3082_/D sky130_fd_sc_hd__nor2_4
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1374_ _2941_/Q _1371_/X _2980_/Q _1372_/X _1373_/X vssd1 vssd1 vccd1 vccd1 _1374_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3044_ _3083_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3044_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2828_ _3101_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2828_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2759_ _2761_/CLK _2759_/D vssd1 vssd1 vccd1 vccd1 _2759_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1992_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__inv_2
XFILLER_159_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2613_ _2700_/Q _2612_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2544_ _2628_/X _2789_/Q _2544_/S vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2475_ _2628_/X _2766_/Q _2475_/S vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1426_ _1426_/A vssd1 vssd1 vccd1 vccd1 _1427_/B sky130_fd_sc_hd__inv_2
XFILLER_29_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1357_ _2861_/Q _1334_/X _1354_/X _1356_/X vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__a211o_1
XFILLER_42_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1288_ _2929_/Q _1269_/X _2968_/Q _1270_/X _1287_/X vssd1 vssd1 vccd1 vccd1 _1288_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3027_ _3105_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3027_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_77_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput570 _2314_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__clkbuf_2
Xoutput581 _2679_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput592 _2689_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _2729_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2260_ vssd1 vssd1 vccd1 vccd1 _2260_/HI _2260_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2191_ _2842_/Q _2157_/X _2186_/X _2190_/X vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__a211o_1
XFILLER_211_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1975_ _2720_/Q _1975_/B vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2527_ _2526_/X _2783_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput309 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 input309/X sky130_fd_sc_hd__buf_1
X_2458_ _2617_/X _2457_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1409_ _3064_/Q _1396_/X _2908_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ _1386_/X _2826_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2389_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _2045_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _2033_/A sky130_fd_sc_hd__or2_2
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1691_ _2788_/Q vssd1 vssd1 vccd1 vccd1 _1691_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2312_ vssd1 vssd1 vccd1 vccd1 _2312_/HI _2312_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2243_ vssd1 vssd1 vccd1 vccd1 _2243_/HI _2243_/LO sky130_fd_sc_hd__conb_1
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2174_ _3074_/Q _2147_/X _2996_/Q _2159_/X vssd1 vssd1 vccd1 vccd1 _2174_/X sky130_fd_sc_hd__a22o_1
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1958_ _1958_/A vssd1 vssd1 vccd1 vccd1 _1959_/B sky130_fd_sc_hd__inv_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1889_ _2695_/Q _1884_/X _2727_/Q _1887_/X vssd1 vssd1 vccd1 vccd1 _2695_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput106 la_data_in[45] vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__buf_1
XPHY_7127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput117 la_data_in[55] vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput128 la_data_in[65] vssd1 vssd1 vccd1 vccd1 _2650_/A0 sky130_fd_sc_hd__clkbuf_2
XPHY_7149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput139 la_data_in[75] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__buf_1
XPHY_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2930_ _3086_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2930_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2861_ _3095_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2861_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_108_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1812_ _1811_/X _1786_/X _1811_/X _1786_/X vssd1 vssd1 vccd1 vccd1 _1812_/Y sky130_fd_sc_hd__a2bb2oi_1
X_2792_ _2792_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2792_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_191_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1743_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1836_/B sky130_fd_sc_hd__buf_2
XFILLER_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1674_ _2765_/Q _1672_/Y _1673_/Y _2789_/Q vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__a22o_1
XFILLER_172_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2226_ vssd1 vssd1 vccd1 vccd1 _2226_/HI _2226_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ _2195_/A vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__buf_1
XPHY_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ _2088_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2553_/S sky130_fd_sc_hd__or2_1
XPHY_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1390_ _2944_/Q _1371_/X _2983_/Q _1372_/X _1389_/X vssd1 vssd1 vccd1 vccd1 _1390_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_122_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3060_ _3099_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3060_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_7480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ _2706_/Q _1947_/B _1948_/A vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__o21a_1
XPHY_6790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2913_ _3108_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2913_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_147_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2844_ _3078_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2844_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_143_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2775_ _2775_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2775_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_199_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1726_ _1724_/Y _2783_/Q _2775_/Q _1725_/Y vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__o22a_1
XFILLER_208_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1657_ _1659_/A _2486_/X vssd1 vssd1 vccd1 vccd1 _2737_/D sky130_fd_sc_hd__and2_1
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1588_ _1533_/B _1582_/B _1533_/B _1582_/B vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2209_ vssd1 vssd1 vccd1 vccd1 _2209_/HI _2209_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2560_ _2721_/Q _2559_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__mux2_1
X_1511_ _1508_/X _1510_/X _1508_/X _1510_/X vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__a2bb2o_1
X_2491_ _2490_/X _2771_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1442_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1443_/B sky130_fd_sc_hd__inv_2
XFILLER_29_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1373_ _3058_/Q _1362_/X _2902_/Q _1363_/X vssd1 vssd1 vccd1 vccd1 _1373_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3112_ _3112_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3112_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_7_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3043_ _3082_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3043_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2827_ _3100_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2827_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_158_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2758_ _2761_/CLK _2758_/D vssd1 vssd1 vccd1 vccd1 _2758_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1709_ _2787_/Q vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2689_ _2722_/CLK _2689_/D vssd1 vssd1 vccd1 vccd1 _2689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1991_ _2725_/Q _1990_/B _1992_/A vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__o21a_1
XFILLER_61_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2612_ _2024_/Y _2700_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2543_ _2542_/X _2788_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2543_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2474_ _2473_/X _2765_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1425_ _1433_/A _1425_/B vssd1 vssd1 vccd1 vccd1 _3074_/D sky130_fd_sc_hd__nor2_4
XFILLER_64_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1356_ _2939_/Q _1337_/X _2978_/Q _1338_/X _1355_/X vssd1 vssd1 vccd1 vccd1 _1356_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1287_ _3046_/Q _1260_/X _2890_/Q _1261_/X vssd1 vssd1 vccd1 vccd1 _1287_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3026_ _3104_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3026_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput560 _2305_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput571 _2664_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput582 _2680_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput593 _2690_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2190_ _2920_/Q _2162_/X _2959_/Q _2164_/X _2189_/X vssd1 vssd1 vccd1 vccd1 _2190_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_211_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1974_ _1974_/A vssd1 vssd1 vccd1 vccd1 _1975_/B sky130_fd_sc_hd__inv_2
XFILLER_109_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2526_ _2628_/X _2783_/Q _2526_/S vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2457_ _2617_/X _2457_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1408_ _3103_/Q _1394_/X _3025_/Q _2109_/A vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__a22o_1
XPHY_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2388_ _1381_/X _2825_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1339_ _3053_/Q _1328_/X _2897_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3009_ _3087_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3009_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput390 _2317_/X vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1690_ _2792_/Q vssd1 vssd1 vccd1 vccd1 _1746_/A sky130_fd_sc_hd__inv_2
XFILLER_32_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2311_ vssd1 vssd1 vccd1 vccd1 _2311_/HI _2311_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2242_ vssd1 vssd1 vccd1 vccd1 _2242_/HI _2242_/LO sky130_fd_sc_hd__conb_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2173_ _2173_/A _2184_/B _2635_/X vssd1 vssd1 vccd1 vccd1 _2800_/D sky130_fd_sc_hd__and3_1
XFILLER_54_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1957_ _2711_/Q _1957_/B vssd1 vssd1 vccd1 vccd1 _1958_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1888_ _2696_/Q _1884_/X _2728_/Q _1887_/X vssd1 vssd1 vccd1 vccd1 _2696_/D sky130_fd_sc_hd__a22o_1
XFILLER_174_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2509_ _2508_/X _2777_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 la_data_in[46] vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__buf_1
XPHY_7128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 la_data_in[56] vssd1 vssd1 vccd1 vccd1 _1478_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput129 la_data_in[66] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__buf_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2860_ _3094_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2860_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ _2767_/Q _2768_/Q _1721_/Y _1666_/Y vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__o22a_1
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2791_ _2791_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2791_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_160_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1742_ _2139_/A _1742_/B vssd1 vssd1 vccd1 vccd1 _2557_/S sky130_fd_sc_hd__nand2_8
XFILLER_102_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1673_ _2765_/Q vssd1 vssd1 vccd1 vccd1 _1673_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2225_ vssd1 vssd1 vccd1 vccd1 _2225_/HI _2225_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2156_ _2156_/A vssd1 vssd1 vccd1 vccd1 _2195_/A sky130_fd_sc_hd__buf_1
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2087_ _2087_/A _2087_/B _2087_/C vssd1 vssd1 vccd1 vccd1 _2550_/S sky130_fd_sc_hd__or3_1
XFILLER_74_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2989_ _3106_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2989_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2010_ _2020_/A _2010_/B vssd1 vssd1 vccd1 vccd1 _2445_/S sky130_fd_sc_hd__and2_4
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _3107_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2912_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2843_ _3077_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2843_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_108_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2774_ _2774_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2774_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_89_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1725_ _2783_/Q vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1656_ _1659_/A _2489_/X vssd1 vssd1 vccd1 vccd1 _2738_/D sky130_fd_sc_hd__and2_1
XFILLER_137_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1587_ _1529_/X _1586_/X _1529_/X _1586_/X vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2208_ vssd1 vssd1 vccd1 vccd1 _2208_/HI _2208_/LO sky130_fd_sc_hd__conb_1
XFILLER_132_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2139_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__buf_1
XFILLER_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1510_ _1443_/B _1509_/X _1443_/B _1509_/X vssd1 vssd1 vccd1 vccd1 _1510_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2490_ _2628_/X _2771_/Q _2490_/S vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1441_ _1445_/A _1441_/B vssd1 vssd1 vccd1 vccd1 _3081_/D sky130_fd_sc_hd__nor2_4
XFILLER_29_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1372_ _2163_/A vssd1 vssd1 vccd1 vccd1 _1372_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3111_ _3111_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3111_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_99_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3042_ _3081_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3042_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput290 la_oenb[96] vssd1 vssd1 vccd1 vccd1 input290/X sky130_fd_sc_hd__buf_1
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2826_ _3099_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2826_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_177_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2757_ _2761_/CLK _2757_/D vssd1 vssd1 vccd1 vccd1 _2757_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1708_ _2791_/Q vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__buf_1
XFILLER_173_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2688_ _2722_/CLK _2688_/D vssd1 vssd1 vccd1 vccd1 _2688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1639_ _1641_/A _2531_/X vssd1 vssd1 vccd1 vccd1 _2752_/D sky130_fd_sc_hd__and2_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1990_ _2725_/Q _1990_/B vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__nand2_1
XFILLER_92_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2611_ _2699_/Q _2610_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2542_ _2541_/X _2788_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2473_ _2472_/X _2765_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1424_ _1424_/A vssd1 vssd1 vccd1 vccd1 _1425_/B sky130_fd_sc_hd__inv_2
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1355_ _3056_/Q _1328_/X _2900_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1355_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1286_ _3085_/Q _1258_/X _3007_/Q _1267_/X vssd1 vssd1 vccd1 vccd1 _1286_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3025_ _3103_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3025_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_23_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2809_ _3082_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2809_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput550 _2296_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput561 _2306_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__clkbuf_2
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput572 _2729_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput583 _2681_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput594 _2691_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1973_ _2719_/Q _1973_/B vssd1 vssd1 vccd1 vccd1 _1974_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2525_ _2524_/X _2782_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2456_ _2615_/X _2455_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1407_ _1417_/A _1611_/B _2392_/X vssd1 vssd1 vccd1 vccd1 _2790_/D sky130_fd_sc_hd__and3_1
XPHY_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2387_ _1375_/X _2824_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1338_ _2199_/A vssd1 vssd1 vccd1 vccd1 _1338_/X sky130_fd_sc_hd__buf_1
XFILLER_211_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1269_ _2198_/A vssd1 vssd1 vccd1 vccd1 _1269_/X sky130_fd_sc_hd__buf_1
XFILLER_186_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3008_ _3086_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3008_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_168_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _2335_/X vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__clkbuf_2
Xoutput391 _2345_/X vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2310_ vssd1 vssd1 vccd1 vccd1 _2310_/HI _2310_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2241_ vssd1 vssd1 vccd1 vccd1 _2241_/HI _2241_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2172_ _2878_/Q _2157_/X _2169_/X _2171_/X vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__a211o_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1956_ _1956_/A vssd1 vssd1 vccd1 vccd1 _1957_/B sky130_fd_sc_hd__inv_2
XFILLER_193_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1887_ _1901_/A vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2508_ _2628_/X _2777_/Q _2508_/S vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 la_data_in[47] vssd1 vssd1 vccd1 vccd1 _1458_/A sky130_fd_sc_hd__buf_1
XFILLER_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2439_ _2600_/X _2439_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2439_/X sky130_fd_sc_hd__mux2_1
Xinput119 la_data_in[57] vssd1 vssd1 vccd1 vccd1 _1481_/A sky130_fd_sc_hd__buf_2
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1810_ _1667_/Y _2770_/Q _2772_/Q _1677_/Y vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__o22a_1
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _2790_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2790_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_106_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1741_ _1688_/X _1740_/X _1688_/X _1740_/X vssd1 vssd1 vccd1 vccd1 _1742_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_106_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1672_ _2789_/Q vssd1 vssd1 vccd1 vccd1 _1672_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2224_ vssd1 vssd1 vccd1 vccd1 _2224_/HI _2224_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2155_ _2173_/A _2184_/B _2633_/X vssd1 vssd1 vccd1 vccd1 _2798_/D sky130_fd_sc_hd__and3_1
XFILLER_61_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2086_ _2086_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2547_/S sky130_fd_sc_hd__or2_1
XFILLER_78_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2988_ _3105_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2988_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_33_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1939_ _2702_/Q _1939_/B vssd1 vssd1 vccd1 vccd1 _1940_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput90 la_data_in[30] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_1
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2911_ _3106_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2911_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_182_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2842_ _3076_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2842_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2773_ _2773_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2773_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_185_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1724_ _2775_/Q vssd1 vssd1 vccd1 vccd1 _1724_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1655_ _1659_/A _2492_/X vssd1 vssd1 vccd1 vccd1 _2739_/D sky130_fd_sc_hd__and2_1
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1586_ _1428_/A _1585_/X _1428_/A _1585_/X vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_113_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2207_ vssd1 vssd1 vccd1 vccd1 _2207_/HI _2207_/LO sky130_fd_sc_hd__conb_1
XFILLER_187_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2138_ _2874_/Q _2102_/X _2135_/X _2137_/X vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__a211o_1
XFILLER_187_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2069_ _2087_/A _2078_/B vssd1 vssd1 vccd1 vccd1 _2505_/S sky130_fd_sc_hd__or2_1
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1440_ _1440_/A vssd1 vssd1 vccd1 vccd1 _1441_/B sky130_fd_sc_hd__inv_2
XFILLER_64_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1371_ _2161_/A vssd1 vssd1 vccd1 vccd1 _1371_/X sky130_fd_sc_hd__buf_1
XFILLER_116_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3110_ _3110_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3110_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3041_ _3080_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3041_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput280 la_oenb[87] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__buf_1
Xinput291 la_oenb[97] vssd1 vssd1 vccd1 vccd1 input291/X sky130_fd_sc_hd__buf_1
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ _3098_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2825_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_192_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2756_ _2761_/CLK _2756_/D vssd1 vssd1 vccd1 vccd1 _2756_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1707_ _2790_/Q _2782_/Q _1705_/Y _1706_/Y vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__o22a_1
X_2687_ _2722_/CLK _2687_/D vssd1 vssd1 vccd1 vccd1 _2687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1638_ _1641_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2753_/D sky130_fd_sc_hd__and2_1
XFILLER_47_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1569_ _1565_/X _1568_/X _1565_/X _1568_/X vssd1 vssd1 vccd1 vccd1 _1569_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2610_ _2022_/X _2699_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2541_ _2628_/X _2788_/Q _2541_/S vssd1 vssd1 vccd1 vccd1 _2541_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2472_ _2628_/X _2765_/Q _2472_/S vssd1 vssd1 vccd1 vccd1 _2472_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1423_ _1494_/A vssd1 vssd1 vccd1 vccd1 _1433_/A sky130_fd_sc_hd__buf_4
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1354_ _3095_/Q _1326_/X _3017_/Q _1335_/X vssd1 vssd1 vccd1 vccd1 _1354_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1285_ _1285_/A _1299_/B _2646_/X vssd1 vssd1 vccd1 vccd1 _2772_/D sky130_fd_sc_hd__and3_1
XFILLER_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3024_ _3102_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3024_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_97_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2808_ _3081_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2808_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_105_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2739_ _2761_/CLK _2739_/D vssd1 vssd1 vccd1 vccd1 _2739_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput540 _2287_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput551 _2297_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput562 _2307_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput573 _2351_/X vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__clkbuf_2
Xoutput584 _2682_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput595 _2692_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1972_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1973_/B sky130_fd_sc_hd__inv_2
XPHY_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2524_ _2523_/X _2782_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2455_ _2615_/X _2455_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1406_ _2192_/A vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2386_ _1366_/X _2823_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1337_ _2198_/A vssd1 vssd1 vccd1 vccd1 _1337_/X sky130_fd_sc_hd__buf_1
XPHY_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1268_ _3082_/Q _1258_/X _3004_/Q _1267_/X vssd1 vssd1 vccd1 vccd1 _1268_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3007_ _3085_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3007_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput370 _2326_/X vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__clkbuf_2
Xoutput381 _2336_/X vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput392 _2346_/X vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2240_ vssd1 vssd1 vccd1 vccd1 _2240_/HI _2240_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2171_ _2956_/Q _2162_/X _2995_/Q _2164_/X _2170_/X vssd1 vssd1 vccd1 vccd1 _2171_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ _2710_/Q _1955_/B vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__nand2_1
XFILLER_202_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1886_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1901_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2507_ _2506_/X _2776_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2507_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput109 la_data_in[48] vssd1 vssd1 vccd1 vccd1 _1460_/A sky130_fd_sc_hd__buf_1
XFILLER_9_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2438_ _2598_/X _2437_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__mux2_1
XPHY_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2369_ _2748_/Q vssd1 vssd1 vccd1 vccd1 _2369_/X sky130_fd_sc_hd__clkbuf_4
XPHY_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _1704_/X _1739_/Y _1704_/X _1739_/Y vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1671_ _1669_/Y _1670_/Y _2776_/Q _2784_/Q vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__a22o_1
XFILLER_176_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2223_ vssd1 vssd1 vccd1 vccd1 _2223_/HI _2223_/LO sky130_fd_sc_hd__conb_1
XFILLER_117_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2154_ _2154_/A vssd1 vssd1 vccd1 vccd1 _2184_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2085_ _2085_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2544_/S sky130_fd_sc_hd__or2_1
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2987_ _3104_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2987_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1938_ _1938_/A vssd1 vssd1 vccd1 vccd1 _1939_/B sky130_fd_sc_hd__inv_2
XFILLER_148_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1869_ _1872_/A _2434_/X vssd1 vssd1 vccd1 vccd1 _2706_/D sky130_fd_sc_hd__and2_1
XFILLER_102_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput80 la_data_in[21] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_1
XFILLER_200_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput91 la_data_in[31] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_1
XFILLER_89_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2910_ _3105_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2910_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_36_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2841_ _3075_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2841_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2772_ _2772_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2772_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1723_ _1721_/Y _2771_/Q _2767_/Q _1722_/Y vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__o22a_1
XFILLER_145_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1654_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1659_/A sky130_fd_sc_hd__buf_1
XFILLER_176_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1585_ _1583_/X _1584_/X _1583_/X _1584_/X vssd1 vssd1 vccd1 vccd1 _1585_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2206_ _2922_/Q _2198_/X _2961_/Q _2199_/X _2205_/X vssd1 vssd1 vccd1 vccd1 _2206_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2137_ _2952_/Q _2114_/X _2991_/Q _2117_/X _2136_/X vssd1 vssd1 vccd1 vccd1 _2137_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2068_ _2087_/C _2081_/B vssd1 vssd1 vccd1 vccd1 _2078_/B sky130_fd_sc_hd__or2_1
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1370_ _3097_/Q _1360_/X _3019_/Q _1369_/X vssd1 vssd1 vccd1 vccd1 _1370_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3040_ _3079_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3040_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput270 la_oenb[78] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__buf_1
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput281 la_oenb[88] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_hd__buf_1
Xinput292 la_oenb[98] vssd1 vssd1 vccd1 vccd1 input292/X sky130_fd_sc_hd__buf_1
XFILLER_23_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2824_ _3097_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2824_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2755_ _2761_/CLK _2755_/D vssd1 vssd1 vccd1 vccd1 _2755_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_30_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1706_ _2782_/Q vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2686_ _2722_/CLK _2686_/D vssd1 vssd1 vccd1 vccd1 _2686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1637_ _1641_/A _2537_/X vssd1 vssd1 vccd1 vccd1 _2754_/D sky130_fd_sc_hd__and2_1
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1568_ _1566_/X _1567_/X _1566_/X _1567_/X vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1499_ _1496_/X _1498_/X _1496_/X _1498_/X vssd1 vssd1 vccd1 vccd1 _1499_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2540_ _2539_/X _2787_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2471_ _2470_/X _2764_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1422_ _1836_/B _1611_/B _2395_/X vssd1 vssd1 vccd1 vccd1 _2793_/D sky130_fd_sc_hd__and3_1
XFILLER_170_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1353_ _1353_/A _1367_/B _2384_/X vssd1 vssd1 vccd1 vccd1 _2782_/D sky130_fd_sc_hd__and3_1
XFILLER_69_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1284_ _2850_/Q _1266_/X _1281_/X _1283_/X vssd1 vssd1 vccd1 vccd1 _1284_/X sky130_fd_sc_hd__a211o_1
XFILLER_62_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3023_ _3101_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3023_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2807_ _3080_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2807_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_121_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2738_ _2761_/CLK _2738_/D vssd1 vssd1 vccd1 vccd1 _2738_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput530 _2223_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__clkbuf_2
X_2669_ _2722_/CLK _2669_/D vssd1 vssd1 vccd1 vccd1 _2669_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput541 _2224_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput552 _2225_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput563 _2226_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput574 _2227_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput585 _2683_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput596 _2693_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1971_ _2718_/Q _1971_/B vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__nand2_1
XPHY_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2523_ _2628_/X _2782_/Q _2523_/S vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2454_ _2613_/X _2453_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1405_ _2868_/Q _2102_/A _1402_/X _1404_/X vssd1 vssd1 vccd1 vccd1 _1405_/X sky130_fd_sc_hd__a211o_1
XFILLER_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2385_ _1357_/X _2822_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1336_ _3092_/Q _1326_/X _3014_/Q _1335_/X vssd1 vssd1 vccd1 vccd1 _1336_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ _2196_/A vssd1 vssd1 vccd1 vccd1 _1267_/X sky130_fd_sc_hd__buf_1
XFILLER_72_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3006_ _3084_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3006_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput371 _2327_/X vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__clkbuf_2
Xoutput382 _2337_/X vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput393 _2347_/X vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2170_ _3073_/Q _2149_/X _2917_/Q _2150_/X vssd1 vssd1 vccd1 vccd1 _2170_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1954_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1955_/B sky130_fd_sc_hd__inv_2
XFILLER_33_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1885_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__inv_2
XFILLER_200_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2506_ _2505_/X _2776_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2437_ _2598_/X _2437_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2368_ _2747_/Q vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1319_ _1319_/A _1333_/B _2652_/X vssd1 vssd1 vccd1 vccd1 _2777_/D sky130_fd_sc_hd__and3_1
XFILLER_61_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2299_ vssd1 vssd1 vccd1 vccd1 _2299_/HI _2299_/LO sky130_fd_sc_hd__conb_1
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1670_ _2784_/Q vssd1 vssd1 vccd1 vccd1 _1670_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2222_ vssd1 vssd1 vccd1 vccd1 _2222_/HI _2222_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2153_ _2876_/Q _2102_/X _2148_/X _2152_/X vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__a211o_1
XFILLER_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2084_ _2084_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2541_/S sky130_fd_sc_hd__or2_1
XFILLER_207_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2986_ _3103_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2986_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1937_ _2701_/Q _2024_/A vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1868_ _1872_/A _2436_/X vssd1 vssd1 vccd1 vccd1 _2707_/D sky130_fd_sc_hd__and2_1
XFILLER_163_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput70 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
XFILLER_102_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput81 la_data_in[22] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_1
Xinput92 la_data_in[32] vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__clkbuf_2
X_1799_ _1746_/X _1798_/X _1746_/X _1798_/X vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_200_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2840_ _3074_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2840_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2771_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2771_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1722_ _2771_/Q vssd1 vssd1 vccd1 vccd1 _1722_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1653_ _1653_/A _2495_/X vssd1 vssd1 vccd1 vccd1 _2740_/D sky130_fd_sc_hd__and2_1
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1584_ _1484_/B _1577_/C _1484_/B _1577_/C vssd1 vssd1 vccd1 vccd1 _1584_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2205_ _3039_/Q _2187_/X _2883_/Q _2188_/X vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__a22o_1
XFILLER_152_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2136_ _3069_/Q _2120_/X _2913_/Q _2124_/X vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2067_ _2086_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2502_/S sky130_fd_sc_hd__or2_1
XFILLER_93_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _3086_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2969_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput260 la_oenb[69] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_hd__buf_1
XFILLER_62_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput271 la_oenb[79] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_hd__buf_1
Xinput282 la_oenb[89] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_hd__buf_1
XFILLER_3_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput293 la_oenb[99] vssd1 vssd1 vccd1 vccd1 input293/X sky130_fd_sc_hd__buf_1
XFILLER_110_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2823_ _3096_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2823_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_207_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2754_ _2761_/CLK _2754_/D vssd1 vssd1 vccd1 vccd1 _2754_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_203_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1705_ _2790_/Q vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2685_ _2722_/CLK _2685_/D vssd1 vssd1 vccd1 vccd1 _2685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1636_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1567_ _1454_/B _1474_/A _1453_/A _1475_/B vssd1 vssd1 vccd1 vccd1 _1567_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1498_ _1472_/A _1497_/X _1472_/A _1497_/X vssd1 vssd1 vccd1 vccd1 _1498_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2119_ _2119_/A vssd1 vssd1 vccd1 vccd1 _2187_/A sky130_fd_sc_hd__buf_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3099_ _3099_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3099_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_58_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2470_ _2469_/X _2764_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1421_ _2871_/Q _2102_/A _1418_/X _1420_/X vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__a211o_1
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1352_ _2860_/Q _1334_/X _1349_/X _1351_/X vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__a211o_1
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1283_ _2928_/Q _1269_/X _2967_/Q _1270_/X _1282_/X vssd1 vssd1 vccd1 vccd1 _1283_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3022_ _3100_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3022_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_62_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2806_ _3079_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2806_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_146_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2737_ _2761_/CLK _2737_/D vssd1 vssd1 vccd1 vccd1 _2737_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2668_ _2722_/CLK _2668_/D vssd1 vssd1 vccd1 vccd1 _2668_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput520 _2268_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput531 _2278_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput542 _2288_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput553 _2298_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__clkbuf_2
X_1619_ _2106_/X _1617_/X _1618_/X _1613_/X vssd1 vssd1 vccd1 vccd1 _1619_/X sky130_fd_sc_hd__o31a_4
Xoutput564 _2308_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2599_ _2014_/X _2709_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__mux2_1
Xoutput575 _2207_/HI vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput586 _2684_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput597 _2694_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1970_ _1970_/A vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__inv_2
XFILLER_72_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2522_ _2521_/X _2781_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2453_ _2613_/X _2453_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1404_ _2946_/Q _2114_/A _2985_/Q _2117_/A _1403_/X vssd1 vssd1 vccd1 vccd1 _1404_/X
+ sky130_fd_sc_hd__a221o_1
X_2384_ _1352_/X _2821_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1335_ _2196_/A vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__buf_1
XFILLER_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_1266_ _2195_/A vssd1 vssd1 vccd1 vccd1 _1266_/X sky130_fd_sc_hd__buf_1
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3005_ _3083_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3005_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_211_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput372 _2328_/X vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput383 _2338_/X vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput394 _2348_/X vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1953_ _2709_/Q _1953_/B vssd1 vssd1 vccd1 vccd1 _1954_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1884_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2505_ _2628_/X _2776_/Q _2505_/S vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2436_ _2596_/X _2435_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2367_ _2746_/Q vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1318_ _2855_/Q _1300_/X _1315_/X _1317_/X vssd1 vssd1 vccd1 vccd1 _1318_/X sky130_fd_sc_hd__a211o_1
XPHY_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2298_ vssd1 vssd1 vccd1 vccd1 _2298_/HI _2298_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1249_ _2845_/Q _2195_/X _1246_/X _1248_/X vssd1 vssd1 vccd1 vccd1 _1249_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_40 _2375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2221_ vssd1 vssd1 vccd1 vccd1 _2221_/HI _2221_/LO sky130_fd_sc_hd__conb_1
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2152_ _2954_/Q _2114_/X _2993_/Q _2117_/X _2151_/X vssd1 vssd1 vccd1 vccd1 _2152_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_66_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2083_ _2087_/B vssd1 vssd1 vccd1 vccd1 _2089_/B sky130_fd_sc_hd__buf_1
XFILLER_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2985_ _3102_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2985_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1936_ _2699_/Q _1936_/B _2700_/Q vssd1 vssd1 vccd1 vccd1 _2024_/A sky130_fd_sc_hd__and3_1
XFILLER_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1867_ _2154_/A vssd1 vssd1 vccd1 vccd1 _1872_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput60 la_data_in[119] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_1
Xinput71 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_1
XFILLER_200_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput82 la_data_in[23] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_1
X_1798_ _1708_/X _1797_/X _1708_/X _1797_/X vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput93 la_data_in[33] vssd1 vssd1 vccd1 vccd1 _1426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2419_ _2580_/X _2419_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _2770_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2770_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ _2767_/Q vssd1 vssd1 vccd1 vccd1 _1721_/Y sky130_fd_sc_hd__inv_2
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1652_ _1653_/A _2498_/X vssd1 vssd1 vccd1 vccd1 _2741_/D sky130_fd_sc_hd__and2_1
XFILLER_12_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1583_ _1464_/B _1563_/C _1464_/B _1563_/C vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2204_ _3078_/Q _2185_/X _3000_/Q _2196_/X vssd1 vssd1 vccd1 vccd1 _2204_/X sky130_fd_sc_hd__a22o_1
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2135_ _3108_/Q _2106_/X _3030_/Q _2109_/X vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2066_ _2081_/B _2085_/A vssd1 vssd1 vccd1 vccd1 _2499_/S sky130_fd_sc_hd__or2_1
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2968_ _3085_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2968_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_210_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1919_ _2673_/Q _1914_/X _2705_/Q _1915_/X vssd1 vssd1 vccd1 vccd1 _2673_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2899_ _3094_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2899_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_198_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput250 la_oenb[5] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__buf_1
XPHY_7271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput261 la_oenb[6] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_hd__buf_1
XPHY_7282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput272 la_oenb[7] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_hd__buf_1
XFILLER_62_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput283 la_oenb[8] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_1
XPHY_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput294 la_oenb[9] vssd1 vssd1 vccd1 vccd1 input294/X sky130_fd_sc_hd__buf_1
XFILLER_209_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2822_ _3095_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2822_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2753_ _2761_/CLK _2753_/D vssd1 vssd1 vccd1 vccd1 _2753_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1704_ _1693_/X _1703_/X _1693_/X _1703_/X vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2684_ _2722_/CLK _2684_/D vssd1 vssd1 vccd1 vccd1 _2684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1635_ _1635_/A _2540_/X vssd1 vssd1 vccd1 vccd1 _2755_/D sky130_fd_sc_hd__and2_1
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1566_ _1456_/B _1482_/B _1455_/A _1481_/A vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1497_ _1447_/A _1454_/B _1448_/B _1453_/A vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2118_ _2398_/S _2118_/B _2118_/C vssd1 vssd1 vccd1 vccd1 _2119_/A sky130_fd_sc_hd__and3_1
X_3098_ _3098_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3098_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_93_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2049_ _2065_/B _2073_/A vssd1 vssd1 vccd1 vccd1 _2076_/A sky130_fd_sc_hd__or2_1
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1420_ _2949_/Q _2114_/A _2988_/Q _2117_/A _1419_/X vssd1 vssd1 vccd1 vccd1 _1420_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1351_ _2938_/Q _1337_/X _2977_/Q _1338_/X _1350_/X vssd1 vssd1 vccd1 vccd1 _1351_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1282_ _3045_/Q _1260_/X _2889_/Q _1261_/X vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3021_ _3099_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3021_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2805_ _3078_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2805_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_160_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2736_ _2761_/CLK _2736_/D vssd1 vssd1 vccd1 vccd1 _2736_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_195_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput510 _2259_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__clkbuf_2
X_2667_ _2722_/CLK _2667_/D vssd1 vssd1 vccd1 vccd1 _2667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput521 _2269_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__clkbuf_2
Xoutput532 _2279_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput543 _2289_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput554 _2299_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__clkbuf_2
X_1618_ _2645_/S _2124_/X _2156_/A vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__or3_4
XFILLER_173_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2598_ _2708_/Q _2597_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__mux2_1
Xoutput565 _2309_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__clkbuf_2
Xoutput576 _2665_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput587 _2666_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput598 _2667_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1549_ _1470_/A _1479_/B _1471_/B _1478_/A vssd1 vssd1 vccd1 vccd1 _1549_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2521_ _2520_/X _2781_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2452_ _2611_/X _2451_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1403_ _3063_/Q _1396_/X _2907_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2383_ _1347_/X _2820_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1334_ _2195_/A vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__buf_1
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1265_ _1285_/A _2203_/B _2643_/X vssd1 vssd1 vccd1 vccd1 _2769_/D sky130_fd_sc_hd__and3_1
XFILLER_84_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3004_ _3082_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3004_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2719_ _2722_/CLK _2719_/D vssd1 vssd1 vccd1 vccd1 _2719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput373 _2329_/X vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__clkbuf_2
Xoutput384 _2339_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput395 _2349_/X vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1952_ _1952_/A vssd1 vssd1 vccd1 vccd1 _1953_/B sky130_fd_sc_hd__inv_2
XFILLER_72_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1883_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_204_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2504_ _2503_/X _2775_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2435_ _2596_/X _2435_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2366_ _2745_/Q vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1317_ _2933_/Q _1303_/X _2972_/Q _1304_/X _1316_/X vssd1 vssd1 vccd1 vccd1 _1317_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2297_ vssd1 vssd1 vccd1 vccd1 _2297_/HI _2297_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1248_ _2923_/Q _2198_/X _2962_/Q _2199_/X _1247_/X vssd1 vssd1 vccd1 vccd1 _1248_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_30 _2365_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_41 _2376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2220_ vssd1 vssd1 vccd1 vccd1 _2220_/HI _2220_/LO sky130_fd_sc_hd__conb_1
XFILLER_191_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2151_ _3071_/Q _2149_/X _2915_/Q _2150_/X vssd1 vssd1 vccd1 vccd1 _2151_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2082_ _2082_/A _2628_/S vssd1 vssd1 vccd1 vccd1 _2087_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2984_ _3101_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2984_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_163_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1935_ _1935_/A vssd1 vssd1 vccd1 vccd1 _1936_/B sky130_fd_sc_hd__inv_2
XFILLER_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1866_ _1866_/A _2438_/X vssd1 vssd1 vccd1 vccd1 _2708_/D sky130_fd_sc_hd__and2_1
XFILLER_175_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_1
Xinput61 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_1
Xinput72 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_1
X_1797_ _1695_/Y _2788_/Q _2799_/Q _1691_/Y vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput83 la_data_in[24] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_1
XFILLER_157_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput94 la_data_in[34] vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2418_ _2578_/X _2417_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2349_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1720_ _1712_/X _1719_/X _1712_/X _1719_/X vssd1 vssd1 vccd1 vccd1 _1720_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1651_ _1653_/A _2501_/X vssd1 vssd1 vccd1 vccd1 _2742_/D sky130_fd_sc_hd__and2_1
XFILLER_86_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1582_ _1582_/A _1582_/B vssd1 vssd1 vccd1 vccd1 _3111_/D sky130_fd_sc_hd__nor2_4
XFILLER_125_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2203_ _2203_/A _2203_/B _2639_/X vssd1 vssd1 vccd1 vccd1 _2765_/D sky130_fd_sc_hd__and3_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2134_ _2134_/A _2146_/B _2630_/X vssd1 vssd1 vccd1 vccd1 _2795_/D sky130_fd_sc_hd__and3_1
XFILLER_110_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2065_ _2065_/A _2065_/B vssd1 vssd1 vccd1 vccd1 _2085_/A sky130_fd_sc_hd__or2_1
XFILLER_93_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2967_ _3084_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2967_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1918_ _2674_/Q _1914_/X _2706_/Q _1915_/X vssd1 vssd1 vccd1 vccd1 _2674_/D sky130_fd_sc_hd__a22o_1
X_2898_ _3093_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2898_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_33_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1849_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput240 la_oenb[50] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_1
XFILLER_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 la_oenb[60] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_hd__buf_1
XFILLER_62_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput262 la_oenb[70] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__buf_1
XFILLER_188_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput273 la_oenb[80] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_hd__buf_1
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput284 la_oenb[90] vssd1 vssd1 vccd1 vccd1 input284/X sky130_fd_sc_hd__buf_1
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput295 wb_clk_i vssd1 vssd1 vccd1 vccd1 _2653_/A1 sky130_fd_sc_hd__buf_4
XFILLER_188_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2821_ _3094_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2821_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2752_ _2761_/CLK _2752_/D vssd1 vssd1 vccd1 vccd1 _2752_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1703_ _1696_/X _1702_/X _1696_/X _1702_/X vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_195_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2683_ _2722_/CLK _2683_/D vssd1 vssd1 vccd1 vccd1 _2683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1634_ _1635_/A _2543_/X vssd1 vssd1 vccd1 vccd1 _2756_/D sky130_fd_sc_hd__and2_1
XFILLER_103_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1565_ _1549_/X _1564_/X _1549_/X _1564_/X vssd1 vssd1 vccd1 vccd1 _1565_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_138_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1496_ _1467_/A _1484_/B _1468_/B _1483_/A vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__a22o_1
XFILLER_80_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2117_ _2117_/A vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__buf_1
XFILLER_110_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3097_ _3097_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3097_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_97_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2048_ _2054_/B vssd1 vssd1 vccd1 vccd1 _2060_/A sky130_fd_sc_hd__buf_1
XFILLER_97_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1350_ _3055_/Q _1328_/X _2899_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1350_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1281_ _3084_/Q _1258_/X _3006_/Q _1267_/X vssd1 vssd1 vccd1 vccd1 _1281_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3020_ _3098_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3020_/Q sky130_fd_sc_hd__dlxtn_1
Xclkbuf_1_0_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _2728_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2804_ _3077_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2804_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_158_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2735_ _2761_/CLK _2735_/D vssd1 vssd1 vccd1 vccd1 _2735_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput500 _2250_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__clkbuf_2
X_2666_ _2722_/CLK _2666_/D vssd1 vssd1 vccd1 vccd1 _2666_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput511 _2260_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput522 _2270_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__clkbuf_2
Xoutput533 _2280_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__clkbuf_2
X_1617_ _1743_/A _1617_/B _2120_/X _2396_/X vssd1 vssd1 vccd1 vccd1 _1617_/X sky130_fd_sc_hd__or4b_4
Xoutput544 _2290_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2597_ _2013_/X _2708_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
Xoutput555 _2300_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput566 _2310_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput577 _2675_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput588 _2685_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__clkbuf_2
X_1548_ _1582_/A _1548_/B vssd1 vssd1 vccd1 vccd1 _3108_/D sky130_fd_sc_hd__nor2_4
XFILLER_173_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput599 _2695_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1479_ _1479_/A _1479_/B vssd1 vssd1 vccd1 vccd1 _3098_/D sky130_fd_sc_hd__nor2_4
XFILLER_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2520_ _2628_/X _2781_/Q _2520_/S vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2451_ _2611_/X _2451_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1402_ _3102_/Q _1394_/X _3024_/Q _2109_/A vssd1 vssd1 vccd1 vccd1 _1402_/X sky130_fd_sc_hd__a22o_1
XFILLER_48_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2382_ _1341_/X _2819_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1333_ _1353_/A _1333_/B _2381_/X vssd1 vssd1 vccd1 vccd1 _2779_/D sky130_fd_sc_hd__and3_1
XFILLER_42_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1264_ _2847_/Q _2195_/X _1259_/X _1263_/X vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__a211o_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XFILLER_209_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3003_ _3081_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3003_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2718_ _2722_/CLK _2718_/D vssd1 vssd1 vccd1 vccd1 _2718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2649_ _1307_/X _2814_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput374 _2330_/X vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput385 _2340_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__clkbuf_2
Xoutput396 _2350_/X vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1951_ _2708_/Q _1951_/B vssd1 vssd1 vccd1 vccd1 _1952_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1882_ _1882_/A _2448_/S vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__nand2_4
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2503_ _2502_/X _2775_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2434_ _2594_/X _2433_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2365_ _2744_/Q vssd1 vssd1 vccd1 vccd1 _2365_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1316_ _3050_/Q _1294_/X _2894_/Q _1295_/X vssd1 vssd1 vccd1 vccd1 _1316_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2296_ vssd1 vssd1 vccd1 vccd1 _2296_/HI _2296_/LO sky130_fd_sc_hd__conb_1
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1247_ _3040_/Q _2187_/X _2884_/Q _2188_/X vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_20 _2735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_31 _2366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_42 _2377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2150_ _2188_/A vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__buf_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2081_ _2081_/A _2081_/B vssd1 vssd1 vccd1 vccd1 _2538_/S sky130_fd_sc_hd__or2_1
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2983_ _3100_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2983_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1934_ _2698_/Q _2697_/Q vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1865_ _1866_/A _2440_/X vssd1 vssd1 vccd1 vccd1 _2709_/D sky130_fd_sc_hd__and2_1
XFILLER_198_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput40 la_data_in[100] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
XFILLER_198_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput51 la_data_in[110] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_1
XFILLER_190_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput62 la_data_in[120] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_1
X_1796_ _2789_/Q _1767_/X _2789_/Q _1767_/X vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput73 la_data_in[15] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_1
Xinput84 la_data_in[25] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_1
XFILLER_196_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput95 la_data_in[35] vssd1 vssd1 vccd1 vccd1 _1430_/A sky130_fd_sc_hd__buf_1
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2417_ _2578_/X _2417_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2348_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2348_/X sky130_fd_sc_hd__clkbuf_1
XPHY_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2279_ vssd1 vssd1 vccd1 vccd1 _2279_/HI _2279_/LO sky130_fd_sc_hd__conb_1
XFILLER_211_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1650_ _1653_/A _2504_/X vssd1 vssd1 vccd1 vccd1 _2743_/D sky130_fd_sc_hd__and2_1
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1581_ _1495_/X _1580_/X _1495_/X _1580_/X vssd1 vssd1 vccd1 vccd1 _1582_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_67_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2202_ _2843_/Q _2195_/X _2197_/X _2201_/X vssd1 vssd1 vccd1 vccd1 _2202_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2133_ _2873_/Q _2102_/X _2130_/X _2132_/X vssd1 vssd1 vccd1 vccd1 _2133_/X sky130_fd_sc_hd__a211o_1
XFILLER_208_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2064_ _2084_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2496_/S sky130_fd_sc_hd__or2_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _3083_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2966_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1917_ _2675_/Q _1914_/X _2707_/Q _1915_/X vssd1 vssd1 vccd1 vccd1 _2675_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2897_ _3092_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2897_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_136_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1848_ _1848_/A _2404_/X vssd1 vssd1 vccd1 vccd1 _2723_/D sky130_fd_sc_hd__and2_1
XFILLER_162_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1779_ _2775_/Q _1778_/Y _1724_/Y _1778_/A vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput230 la_oenb[41] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_1
Xinput241 la_oenb[51] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_1
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput252 la_oenb[61] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__buf_1
XPHY_7273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput263 la_oenb[71] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_hd__buf_1
XPHY_7284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput274 la_oenb[81] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_hd__buf_1
XPHY_7295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput285 la_oenb[91] vssd1 vssd1 vccd1 vccd1 input285/X sky130_fd_sc_hd__buf_1
Xinput296 wb_rst_i vssd1 vssd1 vccd1 vccd1 _2650_/A1 sky130_fd_sc_hd__buf_4
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _3093_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2820_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_143_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ _2761_/CLK _2751_/D vssd1 vssd1 vccd1 vccd1 _2751_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1702_ _2796_/Q _1701_/X _2796_/Q _1701_/X vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_195_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2682_ _2722_/CLK _2682_/D vssd1 vssd1 vccd1 vccd1 _2682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1633_ _1635_/A _2546_/X vssd1 vssd1 vccd1 vccd1 _2757_/D sky130_fd_sc_hd__and2_1
XFILLER_177_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1564_ _1461_/B _1466_/B _1460_/A _1465_/A vssd1 vssd1 vccd1 vccd1 _1564_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1495_ _1487_/A _1491_/A _1488_/B _1492_/B vssd1 vssd1 vccd1 vccd1 _1495_/X sky130_fd_sc_hd__o22a_1
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2116_ _2163_/A vssd1 vssd1 vccd1 vccd1 _2117_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3096_ _3096_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3096_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ _2047_/A _2075_/A vssd1 vssd1 vccd1 vccd1 _2475_/S sky130_fd_sc_hd__or2_1
XFILLER_97_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2949_ _3105_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2949_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1280_ _1285_/A _1299_/B _2645_/X vssd1 vssd1 vccd1 vccd1 _2771_/D sky130_fd_sc_hd__and3_1
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2803_ _3076_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2803_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2734_ _2761_/CLK _2734_/D vssd1 vssd1 vccd1 vccd1 _2734_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_160_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2665_ _2722_/CLK _2665_/D vssd1 vssd1 vccd1 vccd1 _2665_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput501 _2251_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput512 _2261_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__clkbuf_2
Xoutput523 _2271_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput534 _2281_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__clkbuf_2
X_1616_ _1836_/B _1611_/C _2112_/A _1613_/X vssd1 vssd1 vccd1 vccd1 _1616_/X sky130_fd_sc_hd__o31a_4
X_2596_ _2707_/Q _2595_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
Xoutput545 _2291_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__clkbuf_2
Xoutput556 _2301_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__clkbuf_2
Xoutput567 _2311_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput578 _2676_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_2
X_1547_ _1541_/X _1546_/Y _1541_/X _1546_/Y vssd1 vssd1 vccd1 vccd1 _1548_/B sky130_fd_sc_hd__a2bb2o_2
Xoutput589 _2686_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1478_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1479_/B sky130_fd_sc_hd__inv_2
XFILLER_5_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3079_ _3079_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3079_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2450_ _2609_/X _2449_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1401_ _1417_/A _1401_/B _2391_/X vssd1 vssd1 vccd1 vccd1 _2789_/D sky130_fd_sc_hd__and3_1
XFILLER_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2381_ _1332_/X _2818_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2381_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1332_ _2857_/Q _1300_/X _1327_/X _1331_/X vssd1 vssd1 vccd1 vccd1 _1332_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1263_ _2925_/Q _2198_/X _2964_/Q _2199_/X _1262_/X vssd1 vssd1 vccd1 vccd1 _1263_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
XFILLER_211_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3002_ _3080_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3002_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2717_ _2722_/CLK _2717_/D vssd1 vssd1 vccd1 vccd1 _2717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2648_ _1298_/X _2813_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput375 _2331_/X vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2579_ _2003_/X _2715_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput386 _2341_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__clkbuf_2
Xoutput397 _2350_/A vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1950_ _1950_/A vssd1 vssd1 vccd1 vccd1 _1951_/B sky130_fd_sc_hd__inv_2
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1881_ _1881_/A vssd1 vssd1 vccd1 vccd1 _2462_/S sky130_fd_sc_hd__buf_6
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2502_ _2628_/X _2775_/Q _2502_/S vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2433_ _2594_/X _2433_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2364_ _2743_/Q vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1315_ _3089_/Q _1292_/X _3011_/Q _1301_/X vssd1 vssd1 vccd1 vccd1 _1315_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2295_ vssd1 vssd1 vccd1 vccd1 _2295_/HI _2295_/LO sky130_fd_sc_hd__conb_1
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1246_ _3079_/Q _2185_/X _3001_/Q _2196_/X vssd1 vssd1 vccd1 vccd1 _1246_/X sky130_fd_sc_hd__a22o_1
XFILLER_168_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_10 _3109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _2735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_32 _2367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _2664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2080_ _2080_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2535_/S sky130_fd_sc_hd__or2_1
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2982_ _3099_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2982_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1933_ _2557_/S vssd1 vssd1 vccd1 vccd1 _2589_/S sky130_fd_sc_hd__buf_6
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1864_ _1866_/A _2442_/X vssd1 vssd1 vccd1 vccd1 _2710_/D sky130_fd_sc_hd__and2_1
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput30 io_in[36] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput41 la_data_in[101] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 la_data_in[111] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_1
Xinput63 la_data_in[121] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_1
X_1795_ _2062_/A vssd1 vssd1 vccd1 vccd1 _2627_/S sky130_fd_sc_hd__inv_2
XFILLER_190_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput74 la_data_in[16] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_1
Xinput85 la_data_in[26] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_1
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput96 la_data_in[36] vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2416_ _2576_/X _2415_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2347_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2347_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2278_ vssd1 vssd1 vccd1 vccd1 _2278_/HI _2278_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1580_ _1578_/X _1579_/X _1578_/X _1579_/X vssd1 vssd1 vccd1 vccd1 _1580_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2201_ _2921_/Q _2198_/X _2960_/Q _2199_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _2201_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2132_ _2951_/Q _2114_/X _2990_/Q _2117_/X _2131_/X vssd1 vssd1 vccd1 vccd1 _2132_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2063_ _2081_/B vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__buf_1
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2965_ _3082_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2965_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1916_ _2676_/Q _1914_/X _2708_/Q _1915_/X vssd1 vssd1 vccd1 vccd1 _2676_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2896_ _3091_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2896_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1847_ _1848_/A _2406_/X vssd1 vssd1 vccd1 vccd1 _2724_/D sky130_fd_sc_hd__and2_1
XFILLER_11_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1778_ _1778_/A vssd1 vssd1 vccd1 vccd1 _1778_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 la_oenb[32] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_1
XPHY_7241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput231 la_oenb[42] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_1
XFILLER_49_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput242 la_oenb[52] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_1
XPHY_7263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput253 la_oenb[62] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__buf_1
XPHY_7274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput264 la_oenb[72] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_hd__buf_1
XPHY_7285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput275 la_oenb[82] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_hd__buf_1
XPHY_7296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput286 la_oenb[92] vssd1 vssd1 vccd1 vccd1 input286/X sky130_fd_sc_hd__buf_1
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput297 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input297/X sky130_fd_sc_hd__buf_1
XPHY_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2750_ _2761_/CLK _2750_/D vssd1 vssd1 vccd1 vccd1 _2750_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1701_ _2030_/A _1700_/X _2030_/A _1700_/X vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_199_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2681_ _2722_/CLK _2681_/D vssd1 vssd1 vccd1 vccd1 _2681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1632_ _1635_/A _2549_/X vssd1 vssd1 vccd1 vccd1 _2758_/D sky130_fd_sc_hd__and2_1
XFILLER_32_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1563_ _1879_/A _1609_/B _1563_/C vssd1 vssd1 vccd1 vccd1 _3109_/D sky130_fd_sc_hd__and3_2
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1494_ _1494_/A _1494_/B vssd1 vssd1 vccd1 vccd1 _3105_/D sky130_fd_sc_hd__nor2_4
XFILLER_119_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2115_ _2121_/A _2118_/B _2118_/C vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__and3_1
XFILLER_114_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3095_ _3095_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3095_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_167_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2046_ _2061_/B _2073_/A vssd1 vssd1 vccd1 vccd1 _2075_/A sky130_fd_sc_hd__or2_1
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2948_ _3104_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2948_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2879_ _3074_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2879_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2802_ _3075_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2802_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2733_ _2761_/CLK _2733_/D vssd1 vssd1 vccd1 vccd1 _2733_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2664_ _2729_/CLK _2664_/D vssd1 vssd1 vccd1 vccd1 _2664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput502 _2252_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__clkbuf_2
Xoutput513 _2262_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__clkbuf_2
X_1615_ _1836_/B _1611_/C _2122_/A _1613_/X vssd1 vssd1 vccd1 vccd1 _1615_/X sky130_fd_sc_hd__o31a_4
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput524 _2272_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2595_ _2012_/X _2707_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__mux2_1
Xoutput535 _2282_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__clkbuf_2
Xoutput546 _2292_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__clkbuf_2
Xoutput557 _2302_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput568 _2312_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1546_ _1542_/X _1545_/X _1542_/X _1545_/X vssd1 vssd1 vccd1 vccd1 _1546_/Y sky130_fd_sc_hd__o2bb2ai_1
Xoutput579 _2677_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1477_ _1479_/A _1477_/B vssd1 vssd1 vccd1 vccd1 _3097_/D sky130_fd_sc_hd__nor2_4
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3078_ _3078_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3078_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ _2029_/A _2033_/A vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__or2_1
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1400_ _2867_/Q _1368_/X _1395_/X _1399_/X vssd1 vssd1 vccd1 vccd1 _1400_/X sky130_fd_sc_hd__a211o_1
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2380_ _1323_/X _2817_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1331_ _2935_/Q _1303_/X _2974_/Q _1304_/X _1330_/X vssd1 vssd1 vccd1 vccd1 _1331_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1262_ _3042_/Q _1260_/X _2886_/Q _1261_/X vssd1 vssd1 vccd1 vccd1 _1262_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3001_ _3079_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3001_/Q sky130_fd_sc_hd__dlxtn_1
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XFILLER_42_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2716_ _2722_/CLK _2716_/D vssd1 vssd1 vccd1 vccd1 _2716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2647_ _1289_/X _2812_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2578_ _2714_/Q _2577_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__mux2_1
Xoutput376 _2332_/X vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__clkbuf_2
Xoutput387 _2342_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput398 _2208_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__clkbuf_2
X_1529_ _1436_/A _1494_/B _1437_/B _1493_/A vssd1 vssd1 vccd1 vccd1 _1529_/X sky130_fd_sc_hd__a22o_1
XFILLER_141_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1880_ _1880_/A _1880_/B vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__and2_1
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2501_ _2500_/X _2774_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2432_ _2592_/X _2431_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2363_ _2742_/Q vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1314_ _1319_/A _1333_/B _2651_/X vssd1 vssd1 vccd1 vccd1 _2776_/D sky130_fd_sc_hd__and3_1
XFILLER_111_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2294_ vssd1 vssd1 vccd1 vccd1 _2294_/HI _2294_/LO sky130_fd_sc_hd__conb_1
XFILLER_99_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1245_ _2203_/A _2203_/B _2640_/X vssd1 vssd1 vccd1 vccd1 _2766_/D sky130_fd_sc_hd__and3_1
XFILLER_42_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_11 _2730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_22 _2736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 _2368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _2729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2981_ _3098_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2981_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1932_ _2664_/D _1932_/B vssd1 vssd1 vccd1 vccd1 _2507_/S sky130_fd_sc_hd__nor2_8
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1863_ _1866_/A _2444_/X vssd1 vssd1 vccd1 vccd1 _2711_/D sky130_fd_sc_hd__and2_1
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput20 io_in[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
Xinput31 io_in[37] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 la_data_in[102] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
X_1794_ _1832_/A _2082_/A vssd1 vssd1 vccd1 vccd1 _2062_/A sky130_fd_sc_hd__or2_1
Xinput53 la_data_in[112] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_1
Xinput64 la_data_in[122] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
Xinput75 la_data_in[17] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput86 la_data_in[27] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
Xinput97 la_data_in[37] vssd1 vssd1 vccd1 vccd1 _1436_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2415_ _2576_/X _2415_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2415_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2346_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater610 _2645_/S vssd1 vssd1 vccd1 vccd1 _2652_/S sky130_fd_sc_hd__buf_8
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2277_ vssd1 vssd1 vccd1 vccd1 _2277_/HI _2277_/LO sky130_fd_sc_hd__conb_1
XFILLER_211_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2200_ _3038_/Q _2187_/X _2882_/Q _2188_/X vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2131_ _3068_/Q _2120_/X _2912_/Q _2124_/X vssd1 vssd1 vccd1 vccd1 _2131_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2062_ _2062_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2081_/B sky130_fd_sc_hd__or2_2
XFILLER_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2964_ _3081_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2964_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1915_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__buf_1
XFILLER_33_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2895_ _3090_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2895_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1846_ _1848_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _2725_/D sky130_fd_sc_hd__and2_1
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1777_ _1670_/Y _2780_/Q _2784_/Q _1699_/Y vssd1 vssd1 vccd1 vccd1 _1778_/A sky130_fd_sc_hd__o22a_1
XFILLER_144_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2329_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__clkbuf_1
XPHY_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput210 la_oenb[23] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__buf_1
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput221 la_oenb[33] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_1
XFILLER_209_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput232 la_oenb[43] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_1
XPHY_7253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 la_oenb[53] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_1
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput254 la_oenb[63] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__buf_1
XPHY_7275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput265 la_oenb[73] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_hd__buf_1
XPHY_7286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput276 la_oenb[83] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_hd__buf_1
XPHY_7297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput287 la_oenb[93] vssd1 vssd1 vccd1 vccd1 input287/X sky130_fd_sc_hd__buf_1
XPHY_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput298 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input298/X sky130_fd_sc_hd__buf_1
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1700_ _2764_/Q _2780_/Q _1698_/Y _1699_/Y vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__o22a_1
XFILLER_160_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2680_ _2722_/CLK _2680_/D vssd1 vssd1 vccd1 vccd1 _2680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1631_ _1635_/A _2552_/X vssd1 vssd1 vccd1 vccd1 _2759_/D sky130_fd_sc_hd__and2_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1562_ _1555_/X _1561_/Y _1555_/X _1561_/Y vssd1 vssd1 vccd1 vccd1 _1563_/C sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1493_ _1493_/A vssd1 vssd1 vccd1 vccd1 _1494_/B sky130_fd_sc_hd__inv_2
XFILLER_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2114_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__buf_1
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3094_ _3094_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3094_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2045_ _2045_/A _2053_/A _1832_/B vssd1 vssd1 vccd1 vccd1 _2073_/A sky130_fd_sc_hd__or3b_4
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2947_ _3103_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2947_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_108_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2878_ _3112_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2878_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1829_ _1808_/X _1828_/X _1808_/X _1828_/X vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2801_ _3074_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2801_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2732_ _2761_/CLK _2732_/D vssd1 vssd1 vccd1 vccd1 _2732_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2663_ _2659_/X _2660_/X _2661_/X _2662_/X _2053_/B _1834_/A vssd1 vssd1 vccd1 vccd1
+ _2663_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput503 _2253_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__clkbuf_2
X_1614_ _1836_/B _1611_/C _2100_/A _1613_/X vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__o31a_4
XFILLER_173_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput514 _2263_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__clkbuf_2
X_2594_ _2706_/Q _2593_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__mux2_1
Xoutput525 _2273_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__clkbuf_2
Xoutput536 _2283_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput547 _2293_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__clkbuf_2
X_1545_ _1509_/X _1544_/X _1509_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__a2bb2o_1
Xoutput558 _2303_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__clkbuf_2
Xoutput569 _2313_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1476_ _1476_/A vssd1 vssd1 vccd1 vccd1 _1477_/B sky130_fd_sc_hd__inv_2
XFILLER_25_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3077_ _3077_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3077_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2028_ _2704_/Q _1943_/B _1944_/A vssd1 vssd1 vccd1 vccd1 _2028_/X sky130_fd_sc_hd__o21a_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1330_ _3052_/Q _1328_/X _2896_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1330_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1261_ _2188_/A vssd1 vssd1 vccd1 vccd1 _1261_/X sky130_fd_sc_hd__buf_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3000_ _3078_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3000_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_81_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_42_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2715_ _2722_/CLK _2715_/D vssd1 vssd1 vccd1 vccd1 _2715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2646_ _1284_/X _2811_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2577_ _2002_/X _2714_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput377 _2333_/X vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__clkbuf_2
Xoutput388 _2343_/X vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput399 _2318_/X vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__clkbuf_2
X_1528_ _1445_/B _1451_/A _1527_/X _1452_/B vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__o22a_1
XFILLER_29_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1459_ _1468_/A _1459_/B vssd1 vssd1 vccd1 vccd1 _3089_/D sky130_fd_sc_hd__nor2_4
XFILLER_60_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2500_ _2499_/X _2774_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2500_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2431_ _2592_/X _2431_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2431_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2362_ _2741_/Q vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1313_ _2854_/Q _1300_/X _1310_/X _1312_/X vssd1 vssd1 vccd1 vccd1 _1313_/X sky130_fd_sc_hd__a211o_1
X_2293_ vssd1 vssd1 vccd1 vccd1 _2293_/HI _2293_/LO sky130_fd_sc_hd__conb_1
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1244_ _2844_/Q _2195_/X _2204_/X _2206_/X vssd1 vssd1 vccd1 vccd1 _1244_/X sky130_fd_sc_hd__a211o_1
XFILLER_211_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_12 _2740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_23 _2737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_34 _2369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_45 _2728_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2629_ _2127_/X _2833_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2980_ _3097_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2980_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_43_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1931_ _2557_/S vssd1 vssd1 vccd1 vccd1 _2664_/D sky130_fd_sc_hd__clkinv_8
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1862_ _1866_/A _2446_/X vssd1 vssd1 vccd1 vccd1 _2712_/D sky130_fd_sc_hd__and2_1
XFILLER_50_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput21 io_in[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xinput32 io_in[3] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_1
XFILLER_11_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1793_ _1781_/X _1792_/X _1781_/X _1792_/X vssd1 vssd1 vccd1 vccd1 _2082_/A sky130_fd_sc_hd__a2bb2o_1
Xinput43 la_data_in[103] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
XFILLER_174_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput54 la_data_in[113] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_1
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput65 la_data_in[123] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_1
Xinput76 la_data_in[18] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
Xinput87 la_data_in[28] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_1
Xinput98 la_data_in[38] vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2414_ _2574_/X _2413_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2414_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2345_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater611 _2098_/X vssd1 vssd1 vccd1 vccd1 _2645_/S sky130_fd_sc_hd__buf_8
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2276_ vssd1 vssd1 vccd1 vccd1 _2276_/HI _2276_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2130_ _3107_/Q _2106_/X _3029_/Q _2109_/X vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2061_ _2065_/A _2061_/B vssd1 vssd1 vccd1 vccd1 _2084_/A sky130_fd_sc_hd__or2_1
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2963_ _3080_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2963_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_37_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1914_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2894_ _3089_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2894_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1845_ _1848_/A _2410_/X vssd1 vssd1 vccd1 vccd1 _2726_/D sky130_fd_sc_hd__and2_1
XFILLER_102_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1776_ _2033_/A _2626_/S vssd1 vssd1 vccd1 vccd1 _2087_/C sky130_fd_sc_hd__nand2_2
XFILLER_85_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2259_ vssd1 vssd1 vccd1 vccd1 _2259_/HI _2259_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput200 la_oenb[14] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__buf_1
XPHY_7221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput211 la_oenb[24] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_1
XFILLER_42_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput222 la_oenb[34] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_1
XFILLER_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput233 la_oenb[44] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 la_oenb[54] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_1
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput255 la_oenb[64] vssd1 vssd1 vccd1 vccd1 _2653_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput266 la_oenb[74] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_hd__buf_1
XPHY_7287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput277 la_oenb[84] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_hd__buf_1
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput288 la_oenb[94] vssd1 vssd1 vccd1 vccd1 input288/X sky130_fd_sc_hd__buf_1
XPHY_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput299 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input299/X sky130_fd_sc_hd__buf_1
XFILLER_57_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1630_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1635_/A sky130_fd_sc_hd__buf_2
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1561_ _1556_/X _1560_/X _1556_/X _1560_/X vssd1 vssd1 vccd1 vccd1 _1561_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_193_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1492_ _1494_/A _1492_/B vssd1 vssd1 vccd1 vccd1 _3104_/D sky130_fd_sc_hd__nor2_4
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2113_ _2161_/A vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__buf_1
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3093_ _3093_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3093_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _2047_/A _2072_/A vssd1 vssd1 vccd1 vccd1 _2472_/S sky130_fd_sc_hd__or2_1
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2946_ _3102_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2946_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2877_ _3111_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2877_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_178_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1828_ _1671_/X _1827_/X _1671_/X _1827_/X vssd1 vssd1 vccd1 vccd1 _1828_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1759_ _1732_/X _1758_/X _1732_/X _1758_/X vssd1 vssd1 vccd1 vccd1 _1760_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2800_ _2800_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2800_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_53_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2731_ _2761_/CLK _2731_/D vssd1 vssd1 vccd1 vccd1 _2731_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2662_ _1694_/Y _1724_/Y _1787_/Y _1734_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2662_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput504 _2254_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__clkbuf_2
X_1613_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__clkbuf_4
X_2593_ _2011_/X _2706_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__mux2_1
Xoutput515 _2264_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__clkbuf_2
Xoutput526 _2274_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__clkbuf_2
Xoutput537 _2284_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput548 _2294_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__clkbuf_2
X_1544_ _1524_/X _1543_/X _1524_/X _1543_/X vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput559 _2304_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1475_ _1479_/A _1475_/B vssd1 vssd1 vccd1 vccd1 _3096_/D sky130_fd_sc_hd__nor2_4
XFILLER_25_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _3076_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3076_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2027_ _2703_/Q _1941_/B _1942_/A vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__o21a_1
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2929_ _3085_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2929_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1260_ _2187_/A vssd1 vssd1 vccd1 vccd1 _1260_/X sky130_fd_sc_hd__buf_1
XFILLER_133_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_133_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2714_ _2722_/CLK _2714_/D vssd1 vssd1 vccd1 vccd1 _2714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2645_ _1279_/X _2810_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2576_ _2713_/Q _2575_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput378 _2334_/X vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1527_ _1527_/A vssd1 vssd1 vccd1 vccd1 _1527_/X sky130_fd_sc_hd__buf_1
Xoutput389 _2344_/X vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1458_ _1458_/A vssd1 vssd1 vccd1 vccd1 _1459_/B sky130_fd_sc_hd__inv_2
XFILLER_64_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1389_ _3061_/Q _1362_/X _2905_/Q _1363_/X vssd1 vssd1 vccd1 vccd1 _1389_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3059_ _3098_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3059_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2430_ _2590_/X _2429_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2361_ _2740_/Q vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1312_ _2932_/Q _1303_/X _2971_/Q _1304_/X _1311_/X vssd1 vssd1 vccd1 vccd1 _1312_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2292_ vssd1 vssd1 vccd1 vccd1 _2292_/HI _2292_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_13 _2741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_24 _2738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_35 _2370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_46 _2729_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2628_ _2627_/X _2031_/X _2628_/S vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__mux2_8
XFILLER_192_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ _1978_/X _2721_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1930_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2625_/S sky130_fd_sc_hd__inv_4
XFILLER_91_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1861_ _2154_/A vssd1 vssd1 vccd1 vccd1 _1866_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
Xinput22 io_in[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1792_ _1785_/X _1791_/X _1785_/X _1791_/X vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput33 io_in[4] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
XFILLER_11_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput44 la_data_in[104] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
Xinput55 la_data_in[114] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
Xinput66 la_data_in[124] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_1
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput77 la_data_in[19] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_1
XFILLER_85_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput88 la_data_in[29] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_1
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput99 la_data_in[39] vssd1 vssd1 vccd1 vccd1 _1440_/A sky130_fd_sc_hd__buf_1
X_2413_ _2574_/X _2413_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2344_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater612 _2462_/S vssd1 vssd1 vccd1 vccd1 _2448_/S sky130_fd_sc_hd__buf_8
XFILLER_6_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2275_ vssd1 vssd1 vccd1 vccd1 _2275_/HI _2275_/LO sky130_fd_sc_hd__conb_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2060_ _2060_/A _2081_/A vssd1 vssd1 vccd1 vccd1 _2493_/S sky130_fd_sc_hd__or2_1
XFILLER_207_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2962_ _3079_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2962_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1913_ _2677_/Q _1907_/X _2709_/Q _1908_/X vssd1 vssd1 vccd1 vccd1 _2677_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2893_ _3088_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2893_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_206_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1844_ _1848_/A _2412_/X vssd1 vssd1 vccd1 vccd1 _2727_/D sky130_fd_sc_hd__and2_1
XFILLER_50_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1775_ _1775_/A vssd1 vssd1 vccd1 vccd1 _2626_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2327_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2258_ vssd1 vssd1 vccd1 vccd1 _2258_/HI _2258_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2189_ _3037_/Q _2187_/X _2881_/Q _2188_/X vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__a22o_1
XFILLER_57_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput201 la_oenb[15] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__buf_1
XPHY_7222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput212 la_oenb[25] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__buf_1
Xinput223 la_oenb[35] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_1
XPHY_7244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 la_oenb[45] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_1
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_oenb[55] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_1
XPHY_7266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput256 la_oenb[65] vssd1 vssd1 vccd1 vccd1 _2650_/S sky130_fd_sc_hd__clkbuf_2
XPHY_7277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput267 la_oenb[75] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__buf_1
XPHY_7288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput278 la_oenb[85] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_hd__buf_1
XPHY_7299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput289 la_oenb[95] vssd1 vssd1 vccd1 vccd1 input289/X sky130_fd_sc_hd__buf_1
XFILLER_64_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1560_ _1558_/X _1559_/X _1558_/X _1559_/X vssd1 vssd1 vccd1 vccd1 _1560_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_197_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1491_ _1491_/A vssd1 vssd1 vccd1 vccd1 _1492_/B sky130_fd_sc_hd__inv_2
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2112_ _2112_/A vssd1 vssd1 vccd1 vccd1 _2161_/A sky130_fd_sc_hd__inv_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3092_ _3092_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3092_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2043_ _2059_/A _2087_/A vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__or2_1
XFILLER_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2945_ _3101_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2945_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_182_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2876_ _3110_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2876_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1827_ _2792_/Q _1810_/X _2792_/Q _1810_/X vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1758_ _1746_/X _1757_/Y _1746_/X _1757_/Y vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1689_ _2797_/Q vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2730_ _2761_/CLK _2730_/D vssd1 vssd1 vccd1 vccd1 _2730_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_105_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2661_ _1714_/Y _1683_/Y _1669_/Y _1727_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2661_/X sky130_fd_sc_hd__mux4_1
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1612_ _2045_/A _1609_/B _2645_/S _1494_/A vssd1 vssd1 vccd1 vccd1 _1612_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_86_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2592_ _2705_/Q _2591_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__mux2_1
Xoutput505 _2255_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__clkbuf_2
Xoutput516 _2265_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__clkbuf_2
Xoutput527 _2275_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1543_ _1474_/A _1490_/B _1475_/B _1489_/A vssd1 vssd1 vccd1 vccd1 _1543_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput538 _2285_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__clkbuf_2
XFILLER_181_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput549 _2295_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1474_ _1474_/A vssd1 vssd1 vccd1 vccd1 _1475_/B sky130_fd_sc_hd__inv_2
XFILLER_141_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3075_ _3075_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3075_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2026_ _2702_/Q _1939_/B _1940_/A vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2928_ _3084_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2928_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2859_ _3093_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2859_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_168_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2713_ _2722_/CLK _2713_/D vssd1 vssd1 vccd1 vccd1 _2713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2644_ _1273_/X _2809_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2575_ _2000_/X _2713_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput368 _2315_/X vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__clkbuf_2
X_1526_ _1439_/B _1464_/B _1438_/A _1462_/A vssd1 vssd1 vccd1 vccd1 _1526_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput379 _2316_/X vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1457_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1468_/A sky130_fd_sc_hd__buf_4
XFILLER_116_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1388_ _3100_/Q _1360_/X _3022_/Q _1369_/X vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3058_ _3097_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3058_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_43_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2009_ _2705_/Q _1945_/B _1946_/A vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__o21a_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2360_ _2739_/Q vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1311_ _3049_/Q _1294_/X _2893_/Q _1295_/X vssd1 vssd1 vccd1 vccd1 _1311_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2291_ vssd1 vssd1 vccd1 vccd1 _2291_/HI _2291_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_14 _2742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_25 _2739_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 _2371_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2627_ _2658_/X _2663_/X _2627_/S vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2558_ _2557_/X _2793_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1509_ _1463_/A _1481_/A _1462_/A _1482_/B vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__o22a_1
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2489_ _2488_/X _2770_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ _1860_/A _2416_/X vssd1 vssd1 vccd1 vccd1 _2713_/D sky130_fd_sc_hd__and2_1
XFILLER_54_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 io_in[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
X_1791_ _1786_/X _1790_/X _1786_/X _1790_/X vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__o2bb2a_1
Xinput23 io_in[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput34 io_in[5] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput45 la_data_in[105] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
XFILLER_50_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput56 la_data_in[115] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
XFILLER_171_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 la_data_in[125] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_1
XFILLER_89_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput78 la_data_in[1] vssd1 vssd1 vccd1 vccd1 _1609_/B sky130_fd_sc_hd__buf_4
XFILLER_116_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput89 la_data_in[2] vssd1 vssd1 vccd1 vccd1 _2397_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2412_ _2572_/X _2411_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2343_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2274_ vssd1 vssd1 vccd1 vccd1 _2274_/HI _2274_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater613 _2729_/CLK vssd1 vssd1 vccd1 vccd1 _2761_/CLK sky130_fd_sc_hd__buf_12
XFILLER_22_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1989_ _1989_/A vssd1 vssd1 vccd1 vccd1 _1990_/B sky130_fd_sc_hd__inv_2
XFILLER_181_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2961_ _3078_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2961_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_76_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1912_ _2678_/Q _1907_/X _2710_/Q _1908_/X vssd1 vssd1 vccd1 vccd1 _2678_/D sky130_fd_sc_hd__a22o_1
XFILLER_203_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2892_ _3087_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2892_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1843_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1848_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1774_ _1832_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__or2_1
XFILLER_102_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2326_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ vssd1 vssd1 vccd1 vccd1 _2257_/HI _2257_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2188_ _2188_/A vssd1 vssd1 vccd1 vccd1 _2188_/X sky130_fd_sc_hd__buf_1
XFILLER_96_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput202 la_oenb[16] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_1
XFILLER_81_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 la_oenb[26] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_1
XPHY_7234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput224 la_oenb[36] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_1
XPHY_7245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 la_oenb[46] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_1
XPHY_7256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 la_oenb[56] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_1
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput257 la_oenb[66] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__buf_1
XPHY_7278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput268 la_oenb[76] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__buf_1
XPHY_7289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput279 la_oenb[86] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_hd__buf_1
XFILLER_40_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1490_ _1490_/A _1490_/B vssd1 vssd1 vccd1 vccd1 _3103_/D sky130_fd_sc_hd__nor2_4
XFILLER_165_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2111_ _2118_/C _2111_/B vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__or2_2
X_3091_ _3091_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3091_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2042_ _2047_/A _2089_/A vssd1 vssd1 vccd1 vccd1 _2469_/S sky130_fd_sc_hd__or2_1
XFILLER_3_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2944_ _3100_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2944_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_210_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2875_ _3109_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2875_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_198_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1826_ _1753_/A _1825_/A _1753_/Y _1825_/Y vssd1 vssd1 vccd1 vccd1 _1826_/X sky130_fd_sc_hd__o22a_1
XFILLER_198_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1757_ _1751_/X _1756_/X _1751_/X _1756_/X vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_102_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1688_ _1668_/X _1687_/X _1668_/X _1687_/X vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2309_ vssd1 vssd1 vccd1 vccd1 _2309_/HI _2309_/LO sky130_fd_sc_hd__conb_1
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2660_ _1706_/Y _1725_/Y _1699_/Y _1733_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2660_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1611_ _2045_/A _1611_/B _1611_/C vssd1 vssd1 vccd1 vccd1 _1611_/X sky130_fd_sc_hd__and3_4
X_2591_ _2009_/X _2705_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2591_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput506 _2256_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__clkbuf_2
Xoutput517 _2266_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput528 _2276_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1542_ _1493_/A _1502_/Y _1494_/B _1502_/A vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__a22o_1
Xoutput539 _2286_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1473_ _1479_/A _1473_/B vssd1 vssd1 vccd1 vccd1 _3095_/D sky130_fd_sc_hd__nor2_4
XFILLER_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3074_ _3074_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3074_/Q sky130_fd_sc_hd__dlxtn_1
X_2025_ _2701_/Q _2024_/A _1938_/A vssd1 vssd1 vccd1 vccd1 _2025_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ _3083_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2927_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2858_ _3092_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2858_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1809_ _1806_/X _1808_/X _1806_/X _1808_/X vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2789_ _2789_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2789_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2712_ _2722_/CLK _2712_/D vssd1 vssd1 vccd1 vccd1 _2712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2643_ _1264_/X _2808_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2574_ _2728_/Q _2573_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput369 _2325_/X vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1525_ _1522_/X _1524_/X _1522_/X _1524_/X vssd1 vssd1 vccd1 vccd1 _1525_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_82_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1456_ _1456_/A _1456_/B vssd1 vssd1 vccd1 vccd1 _3088_/D sky130_fd_sc_hd__nor2_4
XFILLER_64_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1387_ _1387_/A _1401_/B _2389_/X vssd1 vssd1 vccd1 vccd1 _2787_/D sky130_fd_sc_hd__and3_1
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3057_ _3096_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3057_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2008_ _2720_/Q _1975_/B _1976_/A vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1310_ _3088_/Q _1292_/X _3010_/Q _1301_/X vssd1 vssd1 vccd1 vccd1 _1310_/X sky130_fd_sc_hd__a22o_1
X_2290_ vssd1 vssd1 vccd1 vccd1 _2290_/HI _2290_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_15 _2743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_26 _2354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _2372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2626_ _2625_/X _2029_/X _2626_/S vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2557_ _2556_/X _2793_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1508_ _1506_/X _1507_/X _1506_/X _1507_/X vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2488_ _2487_/X _2770_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1439_ _1445_/A _1439_/B vssd1 vssd1 vccd1 vccd1 _3080_/D sky130_fd_sc_hd__nor2_4
XPHY_6929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3109_ _3109_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3109_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_186_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 io_in[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_141_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ _1788_/X _1789_/X _1788_/X _1789_/X vssd1 vssd1 vccd1 vccd1 _1790_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput24 io_in[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
Xinput35 io_in[6] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput46 la_data_in[106] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
XFILLER_89_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput57 la_data_in[116] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
Xinput68 la_data_in[126] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_1
XFILLER_171_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput79 la_data_in[20] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_1
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2411_ _2572_/X _2411_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2411_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2342_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2273_ vssd1 vssd1 vccd1 vccd1 _2273_/HI _2273_/LO sky130_fd_sc_hd__conb_1
Xrepeater614 _2728_/CLK vssd1 vssd1 vccd1 vccd1 _2722_/CLK sky130_fd_sc_hd__buf_12
XFILLER_26_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1988_ _2724_/Q _1987_/B _1989_/A vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2609_ _2698_/Q _2608_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2960_ _3077_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2960_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1911_ _2679_/Q _1907_/X _2711_/Q _1908_/X vssd1 vssd1 vccd1 vccd1 _2679_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2891_ _3086_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2891_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1842_ _2192_/A vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__buf_2
XFILLER_175_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1773_ _1764_/X _1772_/X _1764_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2325_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2256_ vssd1 vssd1 vccd1 vccd1 _2256_/HI _2256_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2187_ _2187_/A vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__buf_1
XFILLER_187_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput203 la_oenb[17] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__buf_1
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 la_oenb[27] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__buf_1
XPHY_7235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput225 la_oenb[37] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_1
XFILLER_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 la_oenb[47] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_1
XFILLER_44_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput247 la_oenb[57] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__buf_1
XPHY_7268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 la_oenb[67] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__buf_1
XFILLER_44_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput269 la_oenb[77] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__buf_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2110_ _3106_/Q _2106_/X _3028_/Q _2109_/X vssd1 vssd1 vccd1 vccd1 _2110_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3090_ _3090_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3090_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_181_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2041_ _2087_/A _2065_/B vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__or2_1
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2943_ _3099_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2943_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_200_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2874_ _3108_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2874_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1825_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1825_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1756_ _1754_/X _1755_/X _1754_/X _1755_/X vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1687_ _1671_/X _1686_/X _1671_/X _1686_/X vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2308_ vssd1 vssd1 vccd1 vccd1 _2308_/HI _2308_/LO sky130_fd_sc_hd__conb_1
XFILLER_58_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ vssd1 vssd1 vccd1 vccd1 _2239_/HI _2239_/LO sky130_fd_sc_hd__conb_1
XPHY_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1610_ _1617_/B vssd1 vssd1 vccd1 vccd1 _1611_/C sky130_fd_sc_hd__buf_2
XFILLER_103_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2590_ _2720_/Q _2589_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput507 _2257_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__clkbuf_2
Xoutput518 _2267_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1541_ _1536_/X _1540_/X _1536_/X _1540_/X vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput529 _2277_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1472_ _1472_/A vssd1 vssd1 vccd1 vccd1 _1473_/B sky130_fd_sc_hd__inv_2
XFILLER_116_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3073_ _3112_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3073_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2024_ _2024_/A _2024_/B vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2926_ _3082_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2926_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_71_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2857_ _3091_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2857_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1808_ _1722_/Y _2769_/Q _2771_/Q _1807_/Y vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2788_ _2788_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2788_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1739_ _1720_/X _1738_/Y _1720_/X _1738_/Y vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _2722_/CLK _2711_/D vssd1 vssd1 vccd1 vccd1 _2711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2642_ _1255_/X _2807_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2573_ _1999_/X _2728_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1524_ _1431_/B _1523_/X _1431_/B _1523_/X vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1455_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1456_/B sky130_fd_sc_hd__inv_2
XFILLER_206_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1386_ _2865_/Q _1368_/X _1383_/X _1385_/X vssd1 vssd1 vccd1 vccd1 _1386_/X sky130_fd_sc_hd__a211o_1
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3056_ _3095_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3056_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_208_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2007_ _2719_/Q _1973_/B _1974_/A vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__o21a_1
XFILLER_208_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2909_ _3104_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2909_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_16 _2731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_27 _2357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _2373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2625_ _1716_/Y _1713_/Y _2625_/S vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2556_ _2628_/X _2793_/Q _2556_/S vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1507_ _1438_/A _1450_/B _1439_/B _1449_/A vssd1 vssd1 vccd1 vccd1 _1507_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2487_ _2628_/X _2770_/Q _2487_/S vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1438_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1439_/B sky130_fd_sc_hd__inv_2
XPHY_6919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1369_ _2158_/A vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__buf_1
X_3108_ _3108_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3108_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3039_ _3078_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3039_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 io_in[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 io_in[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XFILLER_141_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput36 io_in[7] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XFILLER_200_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput47 la_data_in[107] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_1
XFILLER_176_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput58 la_data_in[117] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
XFILLER_89_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput69 la_data_in[127] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
XFILLER_171_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2410_ _2570_/X _2409_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2410_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2341_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2272_ vssd1 vssd1 vccd1 vccd1 _2272_/HI _2272_/LO sky130_fd_sc_hd__conb_1
XFILLER_65_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater615 _2332_/A vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__buf_8
XFILLER_117_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1987_ _2724_/Q _1987_/B vssd1 vssd1 vccd1 vccd1 _1989_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2608_ _2021_/X _2698_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2539_ _2538_/X _2787_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1910_ _2680_/Q _1907_/X _2712_/Q _1908_/X vssd1 vssd1 vccd1 vccd1 _2680_/D sky130_fd_sc_hd__a22o_1
XFILLER_128_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2890_ _3085_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2890_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _2414_/X _1879_/A vssd1 vssd1 vccd1 vccd1 _2728_/D sky130_fd_sc_hd__and2_1
XFILLER_198_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1772_ _1770_/X _1771_/X _1770_/X _1771_/X vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2324_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2255_ vssd1 vssd1 vccd1 vccd1 _2255_/HI _2255_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2186_ _3076_/Q _2185_/X _2998_/Q _2159_/X vssd1 vssd1 vccd1 vccd1 _2186_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 la_oenb[18] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__buf_1
XFILLER_27_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 la_oenb[28] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_1
XFILLER_62_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput226 la_oenb[38] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__buf_1
XPHY_7247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_oenb[48] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_1
XPHY_7258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 la_oenb[58] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__buf_1
XFILLER_44_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput259 la_oenb[68] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_hd__buf_1
XPHY_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2040_ _2045_/A _2040_/B _1760_/B vssd1 vssd1 vccd1 vccd1 _2065_/B sky130_fd_sc_hd__or3b_4
XFILLER_23_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2942_ _3098_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2942_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2873_ _3107_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2873_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1824_ _2793_/Q _1823_/X _2793_/Q _1823_/X vssd1 vssd1 vccd1 vccd1 _1825_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1755_ _1691_/Y _2794_/Q _2788_/Q _2029_/A vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1686_ _1682_/X _1685_/X _1682_/X _1685_/X vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2307_ vssd1 vssd1 vccd1 vccd1 _2307_/HI _2307_/LO sky130_fd_sc_hd__conb_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ vssd1 vssd1 vccd1 vccd1 _2238_/HI _2238_/LO sky130_fd_sc_hd__conb_1
XFILLER_73_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _3112_/Q _2147_/X _3034_/Q _2159_/X vssd1 vssd1 vccd1 vccd1 _2169_/X sky130_fd_sc_hd__a22o_1
XFILLER_187_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1540_ _1456_/B _1539_/Y _1455_/A _1539_/A vssd1 vssd1 vccd1 vccd1 _1540_/X sky130_fd_sc_hd__o22a_1
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput508 _2221_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput519 _2222_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1471_ _1479_/A _1471_/B vssd1 vssd1 vccd1 vccd1 _3094_/D sky130_fd_sc_hd__nor2_4
XFILLER_190_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ _3111_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3072_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_55_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2023_ _2699_/Q _1936_/B _2700_/Q vssd1 vssd1 vccd1 vccd1 _2024_/B sky130_fd_sc_hd__a21oi_1
XFILLER_97_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2925_ _3081_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2925_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2856_ _3090_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2856_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1807_ _2769_/Q vssd1 vssd1 vccd1 vccd1 _1807_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2787_ _2787_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2787_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_69_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1738_ _1723_/X _1737_/Y _1723_/X _1737_/Y vssd1 vssd1 vccd1 vccd1 _1738_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1669_ _2776_/Q vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2710_ _2722_/CLK _2710_/D vssd1 vssd1 vccd1 vccd1 _2710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2641_ _1249_/X _2806_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2572_ _2727_/Q _2571_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1523_ _1460_/A _1479_/B _1461_/B _1478_/A vssd1 vssd1 vccd1 vccd1 _1523_/X sky130_fd_sc_hd__a22o_1
XFILLER_177_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1454_ _1456_/A _1454_/B vssd1 vssd1 vccd1 vccd1 _3087_/D sky130_fd_sc_hd__nor2_4
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1385_ _2943_/Q _1371_/X _2982_/Q _1372_/X _1384_/X vssd1 vssd1 vccd1 vccd1 _1385_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_206_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3055_ _3094_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3055_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2006_ _2718_/Q _1971_/B _1972_/A vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2908_ _3103_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2908_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_162_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2839_ _3112_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2839_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_121_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_17 _2732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _2363_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_39 _2374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2624_ _1695_/Y _1691_/Y _2625_/S vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2555_ _2554_/X _2792_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1506_ _1424_/A _1427_/B _1425_/B _1426_/A vssd1 vssd1 vccd1 vccd1 _1506_/X sky130_fd_sc_hd__a22o_1
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2486_ _2485_/X _2769_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1437_ _1445_/A _1437_/B vssd1 vssd1 vccd1 vccd1 _3079_/D sky130_fd_sc_hd__nor2_4
XPHY_6909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1368_ _2156_/A vssd1 vssd1 vccd1 vccd1 _1368_/X sky130_fd_sc_hd__buf_1
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3107_ _3107_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3107_/Q sky130_fd_sc_hd__dlxtn_1
X_1299_ _1319_/A _1299_/B _2648_/X vssd1 vssd1 vccd1 vccd1 _2774_/D sky130_fd_sc_hd__and3_1
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3038_ _3077_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3038_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 io_in[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
XFILLER_204_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 io_in[32] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XFILLER_35_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 io_in[8] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_1
XFILLER_141_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 la_data_in[108] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_1
Xinput59 la_data_in[118] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2340_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2271_ vssd1 vssd1 vccd1 vccd1 _2271_/HI _2271_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater616 _2650_/X vssd1 vssd1 vccd1 vccd1 _2332_/A sky130_fd_sc_hd__buf_12
XFILLER_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1986_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1987_/B sky130_fd_sc_hd__inv_2
XFILLER_14_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2607_ _2697_/Q _2019_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__mux2_2
XFILLER_200_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2538_ _2628_/X _2787_/Q _2538_/S vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2469_ _2628_/X _2764_/Q _2469_/S vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _2154_/A vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__clkbuf_4
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1771_ _1672_/Y _1730_/Y _2789_/Q _1730_/A vssd1 vssd1 vccd1 vccd1 _1771_/X sky130_fd_sc_hd__o22a_1
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2323_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2323_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2254_ vssd1 vssd1 vccd1 vccd1 _2254_/HI _2254_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ _2185_/A vssd1 vssd1 vccd1 vccd1 _2185_/X sky130_fd_sc_hd__buf_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1969_ _2717_/Q _1969_/B vssd1 vssd1 vccd1 vccd1 _1970_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput205 la_oenb[19] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__buf_1
XFILLER_66_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput216 la_oenb[29] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_1
XPHY_7237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput227 la_oenb[39] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_1
XFILLER_83_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 la_oenb[49] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_1
XPHY_7259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_oenb[59] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__buf_1
XFILLER_25_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2941_ _3097_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2941_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2872_ _3106_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2872_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1823_ _2796_/Q _1684_/Y _1822_/Y _2763_/Q vssd1 vssd1 vccd1 vccd1 _1823_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1754_ _1668_/X _1753_/Y _1668_/X _1753_/Y vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1685_ _1683_/Y _1684_/Y _2779_/Q _2763_/Q vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__a22o_1
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2306_ vssd1 vssd1 vccd1 vccd1 _2306_/HI _2306_/LO sky130_fd_sc_hd__conb_1
XFILLER_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ vssd1 vssd1 vccd1 vccd1 _2237_/HI _2237_/LO sky130_fd_sc_hd__conb_1
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _2173_/A _2184_/B _2634_/X vssd1 vssd1 vccd1 vccd1 _2799_/D sky130_fd_sc_hd__and3_1
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2099_ _2118_/C _2107_/B vssd1 vssd1 vccd1 vccd1 _2100_/A sky130_fd_sc_hd__or2_2
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput509 _2258_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1470_ _1470_/A vssd1 vssd1 vccd1 vccd1 _1471_/B sky130_fd_sc_hd__inv_2
XFILLER_180_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3071_ _3110_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3071_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_62_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2022_ _2699_/Q _1936_/B _2699_/Q _1936_/B vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2924_ _3080_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2924_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2855_ _3089_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2855_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1806_ _1725_/Y _1778_/A _2783_/Q _1778_/Y vssd1 vssd1 vccd1 vccd1 _1806_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2786_ _2786_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2786_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1737_ _1732_/X _1736_/X _1732_/X _1736_/X vssd1 vssd1 vccd1 vccd1 _1737_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_172_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1668_ _1666_/Y _2772_/Q _2768_/Q _1667_/Y vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__o22a_1
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1599_ _1593_/X _1598_/X _1593_/X _1598_/X vssd1 vssd1 vccd1 vccd1 _1599_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_28_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2640_ _1244_/X _2805_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2571_ _1997_/X _2727_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1522_ _1517_/X _1521_/X _1517_/X _1521_/X vssd1 vssd1 vccd1 vccd1 _1522_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1453_ _1453_/A vssd1 vssd1 vccd1 vccd1 _1454_/B sky130_fd_sc_hd__inv_2
XFILLER_9_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1384_ _3060_/Q _1362_/X _2904_/Q _1363_/X vssd1 vssd1 vccd1 vccd1 _1384_/X sky130_fd_sc_hd__a22o_1
XFILLER_171_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3054_ _3093_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3054_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _2717_/Q _1969_/B _1970_/A vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2907_ _3102_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2907_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_108_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2838_ _3111_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2838_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_191_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2769_ _2769_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2769_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 _2733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_29 _2364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2623_ _1672_/Y _1705_/Y _2625_/S vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2554_ _2553_/X _2792_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1505_ _1502_/Y _1504_/A _1502_/A _1504_/Y vssd1 vssd1 vccd1 vccd1 _1505_/X sky130_fd_sc_hd__o22a_1
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2485_ _2484_/X _2769_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1436_ _1436_/A vssd1 vssd1 vccd1 vccd1 _1437_/B sky130_fd_sc_hd__inv_2
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1367_ _1387_/A _1367_/B _2386_/X vssd1 vssd1 vccd1 vccd1 _2784_/D sky130_fd_sc_hd__and3_1
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3106_ _3106_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3106_/Q sky130_fd_sc_hd__dlxtn_1
X_1298_ _2852_/Q _1266_/X _1293_/X _1297_/X vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__a211o_1
X_3037_ _3076_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3037_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 io_in[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 io_in[33] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 io_in[9] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_1
XFILLER_196_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 la_data_in[109] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_183_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2270_ vssd1 vssd1 vccd1 vccd1 _2270_/HI _2270_/LO sky130_fd_sc_hd__conb_1
XFILLER_191_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater617 _2607_/S vssd1 vssd1 vccd1 vccd1 _2621_/S sky130_fd_sc_hd__buf_8
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1985_ _2723_/Q _1984_/B _1986_/A vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2606_ _2712_/Q _2605_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2537_ _2536_/X _2786_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2468_ _2467_/X _2763_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1419_ _3066_/Q _1396_/X _2910_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1419_/X sky130_fd_sc_hd__a22o_1
XPHY_6729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2399_ _2560_/X _2399_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2399_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _1766_/X _1769_/X _1766_/X _1769_/X vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2322_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2253_ vssd1 vssd1 vccd1 vccd1 _2253_/HI _2253_/LO sky130_fd_sc_hd__conb_1
XFILLER_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2184_ _2203_/A _2184_/B _2637_/X vssd1 vssd1 vccd1 vccd1 _2763_/D sky130_fd_sc_hd__and3_1
XFILLER_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1968_ _1968_/A vssd1 vssd1 vccd1 vccd1 _1969_/B sky130_fd_sc_hd__inv_2
XFILLER_198_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1899_ _2687_/Q _1893_/X _2719_/Q _1894_/X vssd1 vssd1 vccd1 vccd1 _2687_/D sky130_fd_sc_hd__a22o_1
XFILLER_194_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput206 la_oenb[1] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__buf_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 la_oenb[2] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_1
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput228 la_oenb[3] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_1
XPHY_7249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput239 la_oenb[4] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_1
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2940_ _3096_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2940_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_91_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2871_ _3105_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2871_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1822_ _2796_/Q vssd1 vssd1 vccd1 vccd1 _1822_/Y sky130_fd_sc_hd__inv_2
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1753_ _1753_/A vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1684_ _2763_/Q vssd1 vssd1 vccd1 vccd1 _1684_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2305_ vssd1 vssd1 vccd1 vccd1 _2305_/HI _2305_/LO sky130_fd_sc_hd__conb_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2236_ vssd1 vssd1 vccd1 vccd1 _2236_/HI _2236_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2877_/Q _2157_/X _2160_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__a211o_1
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2098_ _2098_/A vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__buf_1
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ _3109_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3070_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_83_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2021_ _2698_/Q _2697_/Q _1935_/A vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2923_ _3079_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2923_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2854_ _3088_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2854_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1805_ _1804_/X _1783_/X _1804_/X _1783_/X vssd1 vssd1 vccd1 vccd1 _1805_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2785_ _2785_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2785_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_15_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1736_ _2769_/Q _1735_/X _2769_/Q _1735_/X vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_201_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1667_ _2772_/Q vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1598_ _1594_/Y _1597_/X _1594_/Y _1597_/X vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2219_ vssd1 vssd1 vccd1 vccd1 _2219_/HI _2219_/LO sky130_fd_sc_hd__conb_1
XFILLER_41_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2570_ _2726_/Q _2569_/X _2607_/S vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1521_ _1518_/X _1520_/X _1518_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_154_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1452_ _1456_/A _1452_/B vssd1 vssd1 vccd1 vccd1 _3086_/D sky130_fd_sc_hd__nor2_4
XFILLER_9_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1383_ _3099_/Q _1360_/X _3021_/Q _1369_/X vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3053_ _3092_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3053_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2004_ _2716_/Q _1967_/B _1968_/A vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__o21a_1
XFILLER_188_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2906_ _3101_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2906_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_162_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2837_ _3110_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2837_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2768_ _2768_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2768_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_191_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1719_ _1715_/X _1718_/X _1715_/X _1718_/X vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__a2bb2o_1
X_2699_ _2722_/CLK _2699_/D vssd1 vssd1 vccd1 vccd1 _2699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_19 _2734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2622_ _1710_/Y _1746_/X _2625_/S vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2553_ _2628_/X _2792_/Q _2553_/S vssd1 vssd1 vccd1 vccd1 _2553_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1504_ _1504_/A vssd1 vssd1 vccd1 vccd1 _1504_/Y sky130_fd_sc_hd__inv_2
X_2484_ _2628_/X _2769_/Q _2484_/S vssd1 vssd1 vccd1 vccd1 _2484_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1435_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__buf_4
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1366_ _2862_/Q _1334_/X _1361_/X _1365_/X vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__a211o_1
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3105_ _3105_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3105_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1297_ _2930_/Q _1269_/X _2969_/Q _1270_/X _1296_/X vssd1 vssd1 vccd1 vccd1 _1297_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3036_ _3075_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3036_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_77_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 io_in[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XFILLER_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 io_in[34] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput39 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater618 input39/X vssd1 vssd1 vccd1 vccd1 _2607_/S sky130_fd_sc_hd__buf_8
XFILLER_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1984_ _2723_/Q _1984_/B vssd1 vssd1 vccd1 vccd1 _1986_/A sky130_fd_sc_hd__nand2_1
XFILLER_198_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2605_ _2017_/X _2712_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2536_ _2535_/X _2786_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2467_ _2466_/X _2763_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1418_ _3105_/Q _1394_/X _3027_/Q _2109_/A vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__a22o_1
XPHY_6719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2398_ _2396_/S _2397_/S _2398_/S vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1349_ _3094_/Q _1326_/X _3016_/Q _1335_/X vssd1 vssd1 vccd1 vccd1 _1349_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3019_ _3097_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3019_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_129_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput490 _2241_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2321_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2321_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2252_ vssd1 vssd1 vccd1 vccd1 _2252_/HI _2252_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2183_ _2841_/Q _2157_/X _2180_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _2183_/X sky130_fd_sc_hd__a211o_1
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1967_ _2716_/Q _1967_/B vssd1 vssd1 vccd1 vccd1 _1968_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1898_ _2688_/Q _1893_/X _2720_/Q _1894_/X vssd1 vssd1 vccd1 vccd1 _2688_/D sky130_fd_sc_hd__a22o_1
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2519_ _2518_/X _2780_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2519_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput207 la_oenb[20] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_1
XPHY_7228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput218 la_oenb[30] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_1
XPHY_7239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput229 la_oenb[40] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_1
XPHY_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2870_ _3104_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2870_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_73_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1821_ _1819_/X _1820_/X _1819_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _1821_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_169_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ _1683_/Y _2787_/Q _2779_/Q _1709_/Y vssd1 vssd1 vccd1 vccd1 _1753_/A sky130_fd_sc_hd__o22a_1
XFILLER_184_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1683_ _2779_/Q vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2304_ vssd1 vssd1 vccd1 vccd1 _2304_/HI _2304_/LO sky130_fd_sc_hd__conb_1
XFILLER_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2235_ vssd1 vssd1 vccd1 vccd1 _2235_/HI _2235_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2166_ _2955_/Q _2162_/X _2994_/Q _2164_/X _2165_/X vssd1 vssd1 vccd1 vccd1 _2166_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2097_ _2121_/A _2118_/B _2107_/A vssd1 vssd1 vccd1 vccd1 _2098_/A sky130_fd_sc_hd__and3_1
XPHY_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2999_ _3077_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _2999_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ _2020_/A _2020_/B vssd1 vssd1 vccd1 vccd1 _2461_/S sky130_fd_sc_hd__and2_4
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2922_ _3078_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2922_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2853_ _3087_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2853_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1804_ _1689_/Y _1678_/Y _2797_/Q _2766_/Q vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__a22o_1
XFILLER_125_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2784_ _2784_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2784_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_89_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1735_ _2781_/Q _2773_/Q _1733_/Y _1734_/Y vssd1 vssd1 vccd1 vccd1 _1735_/X sky130_fd_sc_hd__o22a_1
XFILLER_195_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1666_ _2768_/Q vssd1 vssd1 vccd1 vccd1 _1666_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1597_ _1595_/X _1596_/X _1595_/X _1596_/X vssd1 vssd1 vccd1 vccd1 _1597_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2218_ vssd1 vssd1 vccd1 vccd1 _2218_/HI _2218_/LO sky130_fd_sc_hd__conb_1
XFILLER_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2149_ _2187_/A vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__buf_1
XFILLER_57_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1520_ _1498_/X _1519_/X _1498_/X _1519_/X vssd1 vssd1 vccd1 vccd1 _1520_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1451_ _1451_/A vssd1 vssd1 vccd1 vccd1 _1452_/B sky130_fd_sc_hd__inv_2
XFILLER_9_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1382_ _1387_/A _1401_/B _2388_/X vssd1 vssd1 vccd1 vccd1 _2786_/D sky130_fd_sc_hd__and3_1
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _3091_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3052_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2003_ _2715_/Q _1965_/B _1966_/A vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2905_ _3100_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2905_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2836_ _3109_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2836_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_178_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2767_ _2767_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2767_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1718_ _1716_/Y _2029_/A _2795_/Q _2794_/Q vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2698_ _2722_/CLK _2698_/D vssd1 vssd1 vccd1 vccd1 _2698_/Q sky130_fd_sc_hd__dfxtp_1
X_1649_ _1653_/A _2507_/X vssd1 vssd1 vccd1 vccd1 _2744_/D sky130_fd_sc_hd__and2_1
XFILLER_119_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2621_ _2704_/Q _2620_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2552_ _2551_/X _2791_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__mux2_2
XFILLER_157_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1503_ _1430_/A _1432_/A _1431_/B _1433_/B vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__o22a_1
XFILLER_64_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2483_ _2482_/X _2768_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1434_ _2650_/X vssd1 vssd1 vccd1 vccd1 _1480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1365_ _2940_/Q _1337_/X _2979_/Q _1338_/X _1364_/X vssd1 vssd1 vccd1 vccd1 _1365_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3104_ _3104_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3104_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1296_ _3047_/Q _1294_/X _2891_/Q _1295_/X vssd1 vssd1 vccd1 vccd1 _1296_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _3074_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3035_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_77_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2819_ _3092_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2819_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_in[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 io_in[35] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XFILLER_196_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater608 _2507_/S vssd1 vssd1 vccd1 vccd1 _2558_/S sky130_fd_sc_hd__buf_6
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_register_file.clk_i _2653_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_register_file.clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1983_ _1983_/A vssd1 vssd1 vccd1 vccd1 _1984_/B sky130_fd_sc_hd__inv_2
XFILLER_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2604_ _2711_/Q _2603_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2535_ _2628_/X _2786_/Q _2535_/S vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2466_ _2628_/X _2763_/Q _2466_/S vssd1 vssd1 vccd1 vccd1 _2466_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1417_ _1417_/A _1611_/B _2394_/X vssd1 vssd1 vccd1 vccd1 _2792_/D sky130_fd_sc_hd__and3_1
XFILLER_60_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2397_ _2396_/S _2398_/S _2397_/S vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1348_ _1353_/A _1367_/B _2383_/X vssd1 vssd1 vccd1 vccd1 _2781_/D sky130_fd_sc_hd__and3_1
XFILLER_99_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1279_ _2849_/Q _1266_/X _1276_/X _1278_/X vssd1 vssd1 vccd1 vccd1 _1279_/X sky130_fd_sc_hd__a211o_1
XFILLER_168_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3018_ _3096_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3018_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_77_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput480 _2232_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput491 _2242_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2320_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2251_ vssd1 vssd1 vccd1 vccd1 _2251_/HI _2251_/LO sky130_fd_sc_hd__conb_1
XFILLER_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2182_ _2919_/Q _2162_/X _2958_/Q _2164_/X _2181_/X vssd1 vssd1 vccd1 vccd1 _2182_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1966_ _1966_/A vssd1 vssd1 vccd1 vccd1 _1967_/B sky130_fd_sc_hd__inv_2
XFILLER_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1897_ _2689_/Q _1893_/X _2721_/Q _1894_/X vssd1 vssd1 vccd1 vccd1 _2689_/D sky130_fd_sc_hd__a22o_1
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2518_ _2517_/X _2780_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2518_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput208 la_oenb[21] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_1
XPHY_7229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2449_ _2609_/X _2449_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__mux2_1
Xinput219 la_oenb[31] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_1
XPHY_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ _1708_/X _1763_/X _1708_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1751_ _1679_/X _1750_/Y _1679_/X _1750_/Y vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_15_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1682_ _1674_/X _1681_/X _1674_/X _1681_/X vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2303_ vssd1 vssd1 vccd1 vccd1 _2303_/HI _2303_/LO sky130_fd_sc_hd__conb_1
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2234_ vssd1 vssd1 vccd1 vccd1 _2234_/HI _2234_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2165_ _3072_/Q _2149_/X _2916_/Q _2150_/X vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__a22o_1
XFILLER_94_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2096_ _2118_/C vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__inv_2
XFILLER_39_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2998_ _3076_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _2998_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1949_ _2707_/Q _1949_/B vssd1 vssd1 vccd1 vccd1 _1950_/A sky130_fd_sc_hd__nand2_1
XFILLER_181_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2921_ _3077_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2921_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2852_ _3086_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2852_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1803_ _2627_/S _2628_/S vssd1 vssd1 vccd1 vccd1 _2054_/B sky130_fd_sc_hd__or2_2
XFILLER_160_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2783_ _2783_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2783_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1734_ _2773_/Q vssd1 vssd1 vccd1 vccd1 _1734_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1665_ _1665_/A _2465_/X vssd1 vssd1 vccd1 vccd1 _2730_/D sky130_fd_sc_hd__and2_1
XFILLER_89_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1596_ _1476_/A _1572_/Y _1477_/B _1572_/A vssd1 vssd1 vccd1 vccd1 _1596_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ vssd1 vssd1 vccd1 vccd1 _2217_/HI _2217_/LO sky130_fd_sc_hd__conb_1
XFILLER_132_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2148_ _3110_/Q _2147_/X _3032_/Q _2109_/X vssd1 vssd1 vccd1 vccd1 _2148_/X sky130_fd_sc_hd__a22o_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2079_ _2079_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2532_/S sky130_fd_sc_hd__or2_1
XFILLER_165_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1450_ _1456_/A _1450_/B vssd1 vssd1 vccd1 vccd1 _3085_/D sky130_fd_sc_hd__nor2_4
XFILLER_29_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1381_ _2864_/Q _1368_/X _1378_/X _1380_/X vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3090_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3051_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_7390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2002_ _2714_/Q _1963_/B _1964_/A vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2904_ _3099_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2904_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_182_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2835_ _3108_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2835_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2766_ _2766_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2766_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_145_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1717_ _2794_/Q vssd1 vssd1 vccd1 vccd1 _2029_/A sky130_fd_sc_hd__inv_2
X_2697_ _2729_/CLK _2697_/D vssd1 vssd1 vccd1 vccd1 _2697_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1648_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1653_/A sky130_fd_sc_hd__buf_1
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1579_ _1489_/A _1493_/A _1490_/B _1494_/B vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__o22a_1
XFILLER_154_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2620_ _2028_/X _2704_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2551_ _2550_/X _2791_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1502_ _1502_/A vssd1 vssd1 vccd1 vccd1 _1502_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2482_ _2481_/X _2768_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ _1433_/A _1433_/B vssd1 vssd1 vccd1 vccd1 _3078_/D sky130_fd_sc_hd__nor2_4
XFILLER_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1364_ _3057_/Q _1362_/X _2901_/Q _1363_/X vssd1 vssd1 vccd1 vccd1 _1364_/X sky130_fd_sc_hd__a22o_1
XFILLER_99_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3103_ _3103_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3103_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1295_ _2188_/A vssd1 vssd1 vccd1 vccd1 _1295_/X sky130_fd_sc_hd__buf_1
XFILLER_42_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3034_ _3112_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3034_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2818_ _3091_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2818_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_14_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2749_ _2761_/CLK _2749_/D vssd1 vssd1 vccd1 vccd1 _2749_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_in[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater609 _2589_/S vssd1 vssd1 vccd1 vccd1 _2620_/S sky130_fd_sc_hd__buf_8
XFILLER_78_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1982_ _2722_/Q _1981_/B _1983_/A vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2603_ _2016_/X _2711_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2534_ _2533_/X _2785_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2465_ _2464_/X _2762_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1416_ _2870_/Q _2102_/A _1413_/X _1415_/X vssd1 vssd1 vccd1 vccd1 _1416_/X sky130_fd_sc_hd__a211o_1
XFILLER_64_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2396_ _2111_/B _2107_/B _2396_/S vssd1 vssd1 vccd1 vccd1 _2396_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1347_ _2859_/Q _1334_/X _1344_/X _1346_/X vssd1 vssd1 vccd1 vccd1 _1347_/X sky130_fd_sc_hd__a211o_1
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1278_ _2927_/Q _1269_/X _2966_/Q _1270_/X _1277_/X vssd1 vssd1 vccd1 vccd1 _1278_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_211_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3017_ _3095_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3017_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput470 _2372_/X vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput481 _2233_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput492 _2243_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2250_ vssd1 vssd1 vccd1 vccd1 _2250_/HI _2250_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2181_ _3036_/Q _2149_/X _2880_/Q _2150_/X vssd1 vssd1 vccd1 vccd1 _2181_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1965_ _2715_/Q _1965_/B vssd1 vssd1 vccd1 vccd1 _1966_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1896_ _2690_/Q _1893_/X _2722_/Q _1894_/X vssd1 vssd1 vccd1 vccd1 _2690_/D sky130_fd_sc_hd__a22o_1
XFILLER_174_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2517_ _2628_/X _2780_/Q _2517_/S vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2448_ _2607_/X _2447_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2448_/X sky130_fd_sc_hd__mux2_1
Xinput209 la_oenb[22] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__buf_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ _2758_/Q vssd1 vssd1 vccd1 vccd1 _2379_/X sky130_fd_sc_hd__buf_2
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1750_ _1747_/X _1749_/X _1747_/X _1749_/X vssd1 vssd1 vccd1 vccd1 _1750_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_89_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1681_ _1675_/X _1680_/X _1675_/X _1680_/X vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_184_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2302_ vssd1 vssd1 vccd1 vccd1 _2302_/HI _2302_/LO sky130_fd_sc_hd__conb_1
XFILLER_119_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2233_ vssd1 vssd1 vccd1 vccd1 _2233_/HI _2233_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2164_ _2199_/A vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__buf_1
X_2095_ _2396_/S vssd1 vssd1 vccd1 vccd1 _2118_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2997_ _3075_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _2997_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1948_ _1948_/A vssd1 vssd1 vccd1 vccd1 _1949_/B sky130_fd_sc_hd__inv_2
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1879_ _1879_/A _2448_/X vssd1 vssd1 vccd1 vccd1 _2697_/D sky130_fd_sc_hd__and2_1
XFILLER_11_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2920_ _3076_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2920_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2851_ _3085_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2851_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_182_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1802_ _1802_/A vssd1 vssd1 vccd1 vccd1 _2628_/S sky130_fd_sc_hd__buf_1
XFILLER_54_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2782_ _2782_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2782_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1733_ _2781_/Q vssd1 vssd1 vccd1 vccd1 _1733_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1664_ _1665_/A _2468_/X vssd1 vssd1 vccd1 vccd1 _2731_/D sky130_fd_sc_hd__and2_1
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1595_ _1468_/B _1487_/A _1467_/A _1488_/B vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2216_ vssd1 vssd1 vccd1 vccd1 _2216_/HI _2216_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2147_ _2185_/A vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__buf_1
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2078_ _2078_/A _2078_/B vssd1 vssd1 vccd1 vccd1 _2529_/S sky130_fd_sc_hd__or2_1
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1380_ _2942_/Q _1371_/X _2981_/Q _1372_/X _1379_/X vssd1 vssd1 vccd1 vccd1 _1380_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3050_ _3089_/D _1621_/X vssd1 vssd1 vccd1 vccd1 _3050_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_7380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2001_ _2020_/A _2001_/B vssd1 vssd1 vccd1 vccd1 _2429_/S sky130_fd_sc_hd__and2_4
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2903_ _3098_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2903_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2834_ _3107_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2834_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2765_ _2765_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2765_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1716_ _2795_/Q vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2696_ _2728_/CLK _2696_/D vssd1 vssd1 vccd1 vccd1 _2696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1647_ _1647_/A _2510_/X vssd1 vssd1 vccd1 vccd1 _2745_/D sky130_fd_sc_hd__and2_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1578_ _1484_/B _1486_/B _1483_/A _1485_/A vssd1 vssd1 vccd1 vccd1 _1578_/X sky130_fd_sc_hd__a22o_1
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2550_ _2628_/X _2791_/Q _2550_/S vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1501_ _1459_/B _1476_/A _1458_/A _1477_/B vssd1 vssd1 vccd1 vccd1 _1502_/A sky130_fd_sc_hd__o22a_1
XFILLER_157_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2481_ _2628_/X _2768_/Q _2481_/S vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1432_ _1432_/A vssd1 vssd1 vccd1 vccd1 _1433_/B sky130_fd_sc_hd__inv_2
XFILLER_64_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1363_ _2123_/A vssd1 vssd1 vccd1 vccd1 _1363_/X sky130_fd_sc_hd__buf_1
XFILLER_64_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3102_ _3102_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3102_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1294_ _2187_/A vssd1 vssd1 vccd1 vccd1 _1294_/X sky130_fd_sc_hd__buf_1
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3033_ _3111_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3033_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2817_ _3090_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2817_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_53_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2748_ _2761_/CLK _2748_/D vssd1 vssd1 vccd1 vccd1 _2748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2679_ _2722_/CLK _2679_/D vssd1 vssd1 vccd1 vccd1 _2679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1981_ _2722_/Q _1981_/B vssd1 vssd1 vccd1 vccd1 _1983_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2602_ _2710_/Q _2601_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2533_ _2532_/X _2785_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2464_ _2463_/X _2762_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1415_ _2948_/Q _2114_/A _2987_/Q _2117_/A _1414_/X vssd1 vssd1 vccd1 vccd1 _1415_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2395_ _1421_/X _2832_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2395_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1346_ _2937_/Q _1337_/X _2976_/Q _1338_/X _1345_/X vssd1 vssd1 vccd1 vccd1 _1346_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_151_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1277_ _3044_/Q _1260_/X _2888_/Q _1261_/X vssd1 vssd1 vccd1 vccd1 _1277_/X sky130_fd_sc_hd__a22o_1
XFILLER_211_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3016_ _3094_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3016_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput460 _2363_/X vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput471 _2373_/X vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__clkbuf_2
Xoutput482 _2234_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput493 _2244_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2180_ _3075_/Q _2147_/X _2997_/Q _2159_/X vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__a22o_1
XFILLER_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1964_ _1964_/A vssd1 vssd1 vccd1 vccd1 _1965_/B sky130_fd_sc_hd__inv_2
XFILLER_202_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1895_ _2691_/Q _1893_/X _2723_/Q _1894_/X vssd1 vssd1 vccd1 vccd1 _2691_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2516_ _2515_/X _2779_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2516_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2447_ _2607_/X _2447_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2447_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2378_ _2757_/Q vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__buf_2
XFILLER_97_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ _2123_/A vssd1 vssd1 vccd1 vccd1 _1329_/X sky130_fd_sc_hd__buf_1
XPHY_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1680_ _1676_/Y _1679_/X _1676_/Y _1679_/X vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2301_ vssd1 vssd1 vccd1 vccd1 _2301_/HI _2301_/LO sky130_fd_sc_hd__conb_1
XFILLER_48_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2232_ vssd1 vssd1 vccd1 vccd1 _2232_/HI _2232_/LO sky130_fd_sc_hd__conb_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2163_ _2163_/A vssd1 vssd1 vccd1 vccd1 _2199_/A sky130_fd_sc_hd__buf_1
XFILLER_26_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2094_/A vssd1 vssd1 vccd1 vccd1 _2107_/B sky130_fd_sc_hd__buf_1
XFILLER_78_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2996_ _3074_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _2996_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_206_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1947_ _2706_/Q _1947_/B vssd1 vssd1 vccd1 vccd1 _1948_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _1878_/A _2450_/X vssd1 vssd1 vccd1 vccd1 _2698_/D sky130_fd_sc_hd__and2_1
XFILLER_15_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2850_ _3084_/D _1614_/X vssd1 vssd1 vccd1 vccd1 _2850_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1801_ _2139_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _1802_/A sky130_fd_sc_hd__and2_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _2781_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2781_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1732_ _1730_/A _1731_/A _1730_/Y _1731_/Y vssd1 vssd1 vccd1 vccd1 _1732_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1663_ _1665_/A _2471_/X vssd1 vssd1 vccd1 vccd1 _2732_/D sky130_fd_sc_hd__and2_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1594_ _1516_/A _1537_/X _1516_/A _1537_/X vssd1 vssd1 vccd1 vccd1 _1594_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_193_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2215_ vssd1 vssd1 vccd1 vccd1 _2215_/HI _2215_/LO sky130_fd_sc_hd__conb_1
XFILLER_113_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2146_ _2173_/A _2146_/B _2632_/X vssd1 vssd1 vccd1 vccd1 _2797_/D sky130_fd_sc_hd__and3_1
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2077_ _2077_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2526_/S sky130_fd_sc_hd__or2_1
XFILLER_179_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2979_ _3096_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2979_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput360 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 _2431_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2000_ _2713_/Q _1961_/B _1962_/A vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2902_ _3097_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2902_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_71_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2833_ _3106_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2833_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2764_ _2764_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2764_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_145_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1715_ _1713_/Y _2778_/Q _2762_/Q _1714_/Y vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__o22a_1
XFILLER_145_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2695_ _2729_/CLK _2695_/D vssd1 vssd1 vccd1 vccd1 _2695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1646_ _1647_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2746_/D sky130_fd_sc_hd__and2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1577_ _2146_/B _1609_/B _1577_/C vssd1 vssd1 vccd1 vccd1 _3110_/D sky130_fd_sc_hd__and3_2
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2129_ _2134_/A _2146_/B _2629_/X vssd1 vssd1 vccd1 vccd1 _2794_/D sky130_fd_sc_hd__and3_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1500_ _1495_/X _1499_/X _1495_/X _1499_/X vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2480_ _2479_/X _2767_/Q _2507_/S vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1431_ _1433_/A _1431_/B vssd1 vssd1 vccd1 vccd1 _3077_/D sky130_fd_sc_hd__nor2_4
XFILLER_68_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1362_ _2119_/A vssd1 vssd1 vccd1 vccd1 _1362_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3101_ _3101_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3101_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_116_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1293_ _3086_/Q _1292_/X _3008_/Q _1267_/X vssd1 vssd1 vccd1 vccd1 _1293_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3032_ _3110_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3032_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_168_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput190 la_oenb[120] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__buf_1
XFILLER_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2816_ _3089_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2816_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2747_ _2761_/CLK _2747_/D vssd1 vssd1 vccd1 vccd1 _2747_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2678_ _2722_/CLK _2678_/D vssd1 vssd1 vccd1 vccd1 _2678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1629_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1980_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1981_/B sky130_fd_sc_hd__inv_2
XPHY_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2601_ _2015_/X _2710_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2532_ _2628_/X _2785_/Q _2532_/S vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2463_ _2628_/X _2762_/Q _2463_/S vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1414_ _3065_/Q _1396_/X _2909_/Q _1397_/X vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2394_ _1416_/X _2831_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2394_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1345_ _3054_/Q _1328_/X _2898_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1345_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1276_ _3083_/Q _1258_/X _3005_/Q _1267_/X vssd1 vssd1 vccd1 vccd1 _1276_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3015_ _3093_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3015_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_149_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput450 _2354_/X vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput461 _2364_/X vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput472 _2374_/X vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput483 _2235_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput494 _2245_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1963_ _2714_/Q _1963_/B vssd1 vssd1 vccd1 vccd1 _1964_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1894_ _1901_/A vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2515_ _2514_/X _2779_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2515_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2446_ _2606_/X _2445_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2377_ _2756_/Q vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__buf_2
XFILLER_190_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1328_ _2119_/A vssd1 vssd1 vccd1 vccd1 _1328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1259_ _3081_/Q _1258_/X _3003_/Q _2196_/X vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__a22o_1
XFILLER_209_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2300_ vssd1 vssd1 vccd1 vccd1 _2300_/HI _2300_/LO sky130_fd_sc_hd__conb_1
XFILLER_135_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2231_ vssd1 vssd1 vccd1 vccd1 _2231_/HI _2231_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2162_ _2198_/A vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__buf_1
XFILLER_120_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2093_ _2398_/S _2118_/B vssd1 vssd1 vccd1 vccd1 _2094_/A sky130_fd_sc_hd__or2_1
XFILLER_207_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2995_ _3112_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2995_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1946_ _1946_/A vssd1 vssd1 vccd1 vccd1 _1947_/B sky130_fd_sc_hd__inv_2
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1877_ _1878_/A _2452_/X vssd1 vssd1 vccd1 vccd1 _2699_/D sky130_fd_sc_hd__and2_1
XFILLER_50_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2429_ _2590_/X _2429_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2429_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ _1796_/X _1799_/X _1796_/X _1799_/X vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__a2bb2o_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2780_ _2780_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2780_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_180_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1731_ _1731_/A vssd1 vssd1 vccd1 vccd1 _1731_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1662_ _1665_/A _2474_/X vssd1 vssd1 vccd1 vccd1 _2733_/D sky130_fd_sc_hd__and2_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1593_ _1486_/B _1489_/A _1485_/A _1490_/B vssd1 vssd1 vccd1 vccd1 _1593_/X sky130_fd_sc_hd__o22a_1
XFILLER_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2214_ vssd1 vssd1 vccd1 vccd1 _2214_/HI _2214_/LO sky130_fd_sc_hd__conb_1
XFILLER_117_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2145_ _2875_/Q _2102_/X _2142_/X _2144_/X vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__a211o_1
XFILLER_67_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2076_ _2076_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2523_/S sky130_fd_sc_hd__or2_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2978_ _3095_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2978_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1929_ _2665_/Q _1900_/A _2697_/Q _1901_/A vssd1 vssd1 vccd1 vccd1 _2665_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput350 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 _2407_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput361 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 _2433_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2901_ _3096_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2901_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_189_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2832_ _3105_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2832_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_207_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2763_ _2763_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2763_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1714_ _2778_/Q vssd1 vssd1 vccd1 vccd1 _1714_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2694_ _2729_/CLK _2694_/D vssd1 vssd1 vccd1 vccd1 _2694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1645_ _1647_/A _2516_/X vssd1 vssd1 vccd1 vccd1 _2747_/D sky130_fd_sc_hd__and2_1
XFILLER_160_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1576_ _1569_/X _1575_/X _1569_/X _1575_/X vssd1 vssd1 vccd1 vccd1 _1577_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _2192_/A vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2059_/A _2078_/A vssd1 vssd1 vccd1 vccd1 _2081_/A sky130_fd_sc_hd__or2_1
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1430_ _1430_/A vssd1 vssd1 vccd1 vccd1 _1431_/B sky130_fd_sc_hd__inv_2
XFILLER_99_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1361_ _3096_/Q _1360_/X _3018_/Q _1335_/X vssd1 vssd1 vccd1 vccd1 _1361_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3100_ _3100_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3100_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_1_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1292_ _2185_/A vssd1 vssd1 vccd1 vccd1 _1292_/X sky130_fd_sc_hd__buf_1
XFILLER_209_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3031_ _3109_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3031_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_62_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 la_oenb[111] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_hd__buf_1
XFILLER_3_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput191 la_oenb[121] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__buf_1
XFILLER_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2815_ _3088_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2815_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_140_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2746_ _2761_/CLK _2746_/D vssd1 vssd1 vccd1 vccd1 _2746_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2677_ _2722_/CLK _2677_/D vssd1 vssd1 vccd1 vccd1 _2677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1628_ _2139_/A vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1559_ _1438_/A _1482_/B _1439_/B _1481_/A vssd1 vssd1 vccd1 vccd1 _1559_/X sky130_fd_sc_hd__a22o_1
XFILLER_47_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2600_ _2709_/Q _2599_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2531_ _2530_/X _2784_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2462_ _2621_/X _2461_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1413_ _3104_/Q _1394_/X _3026_/Q _2109_/A vssd1 vssd1 vccd1 vccd1 _1413_/X sky130_fd_sc_hd__a22o_1
X_2393_ _1411_/X _2830_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1344_ _3093_/Q _1326_/X _3015_/Q _1335_/X vssd1 vssd1 vccd1 vccd1 _1344_/X sky130_fd_sc_hd__a22o_1
XFILLER_69_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1275_ _1285_/A _1299_/B _2644_/X vssd1 vssd1 vccd1 vccd1 _2770_/D sky130_fd_sc_hd__and3_1
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3014_ _3092_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3014_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_3_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2729_ _2729_/CLK _2729_/D vssd1 vssd1 vccd1 vccd1 _2729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput440 _2736_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput451 _2355_/X vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__clkbuf_2
Xoutput462 _2365_/X vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput473 _2375_/X vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput484 _2236_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput495 _2246_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _1962_/A vssd1 vssd1 vccd1 vccd1 _1963_/B sky130_fd_sc_hd__inv_2
XFILLER_37_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1893_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2514_ _2628_/X _2779_/Q _2514_/S vssd1 vssd1 vccd1 vccd1 _2514_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2445_ _2606_/X _2445_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2376_ _2755_/Q vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1327_ _3091_/Q _1326_/X _3013_/Q _1301_/X vssd1 vssd1 vccd1 vccd1 _1327_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1258_ _2185_/A vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__buf_1
XFILLER_209_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ vssd1 vssd1 vccd1 vccd1 _2230_/HI _2230_/LO sky130_fd_sc_hd__conb_1
XFILLER_117_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2161_ _2161_/A vssd1 vssd1 vccd1 vccd1 _2198_/A sky130_fd_sc_hd__buf_1
XFILLER_117_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2092_ _2121_/A _2118_/B vssd1 vssd1 vccd1 vccd1 _2111_/B sky130_fd_sc_hd__or2_1
XFILLER_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2994_ _3111_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2994_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_203_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1945_ _2705_/Q _1945_/B vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__nand2_1
XFILLER_206_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1876_ _1878_/A _2454_/X vssd1 vssd1 vccd1 vccd1 _2700_/D sky130_fd_sc_hd__and2_1
XFILLER_159_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2428_ _2588_/X _2427_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2359_ _2738_/Q vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ _1730_/A vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1661_ _1665_/A _2477_/X vssd1 vssd1 vccd1 vccd1 _2734_/D sky130_fd_sc_hd__and2_1
XFILLER_125_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1592_ _1491_/A _1504_/Y _1492_/B _1504_/A vssd1 vssd1 vccd1 vccd1 _1592_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2213_ vssd1 vssd1 vccd1 vccd1 _2213_/HI _2213_/LO sky130_fd_sc_hd__conb_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2144_ _2953_/Q _2114_/X _2992_/Q _2117_/X _2143_/X vssd1 vssd1 vccd1 vccd1 _2144_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2075_ _2075_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2520_/S sky130_fd_sc_hd__or2_1
XFILLER_187_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2977_ _3094_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2977_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1928_ _2666_/Q _1900_/A _2698_/Q _1901_/A vssd1 vssd1 vccd1 vccd1 _2666_/D sky130_fd_sc_hd__a22o_1
XFILLER_175_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1859_ _1860_/A _2418_/X vssd1 vssd1 vccd1 vccd1 _2714_/D sky130_fd_sc_hd__and2_1
XFILLER_190_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput340 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 _2421_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput351 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 _2409_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput362 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _2020_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2900_ _3095_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2900_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_127_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2831_ _3104_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2831_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_34_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2762_ _2762_/D _1611_/X vssd1 vssd1 vccd1 vccd1 _2762_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_157_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1713_ _2762_/Q vssd1 vssd1 vccd1 vccd1 _1713_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2693_ _2728_/CLK _2693_/D vssd1 vssd1 vccd1 vccd1 _2693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_0 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1644_ _1647_/A _2519_/X vssd1 vssd1 vccd1 vccd1 _2748_/D sky130_fd_sc_hd__and2_1
XFILLER_138_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1575_ _1570_/X _1574_/X _1570_/X _1574_/X vssd1 vssd1 vccd1 vccd1 _1575_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2127_ _2872_/Q _2102_/X _2110_/X _2126_/X vssd1 vssd1 vccd1 vccd1 _2127_/X sky130_fd_sc_hd__a211o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2058_ _2060_/A _2080_/A vssd1 vssd1 vccd1 vccd1 _2490_/S sky130_fd_sc_hd__or2_1
XFILLER_93_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1360_ _2105_/A vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__buf_1
XFILLER_155_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1291_ _1319_/A _1299_/B _2647_/X vssd1 vssd1 vccd1 vccd1 _2773_/D sky130_fd_sc_hd__and3_1
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3030_ _3108_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3030_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_114_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput170 la_oenb[102] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__buf_1
XFILLER_62_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput181 la_oenb[112] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_hd__buf_1
XFILLER_114_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput192 la_oenb[122] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__buf_1
XFILLER_149_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2814_ _3087_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2814_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2745_ _2761_/CLK _2745_/D vssd1 vssd1 vccd1 vccd1 _2745_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2676_ _2722_/CLK _2676_/D vssd1 vssd1 vccd1 vccd1 _2676_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput600 _2696_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1627_ _2555_/X _2134_/A vssd1 vssd1 vccd1 vccd1 _2760_/D sky130_fd_sc_hd__and2_2
XFILLER_86_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1558_ _1474_/A _1557_/X _1474_/A _1557_/X vssd1 vssd1 vccd1 vccd1 _1558_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1489_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1490_/B sky130_fd_sc_hd__inv_2
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2530_ _2529_/X _2784_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2461_ _2621_/X _2461_/A1 _2461_/S vssd1 vssd1 vccd1 vccd1 _2461_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1412_ _1417_/A _1611_/B _2393_/X vssd1 vssd1 vccd1 vccd1 _2791_/D sky130_fd_sc_hd__and3_1
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2392_ _1405_/X _2829_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1343_ _1353_/A _1367_/B _2382_/X vssd1 vssd1 vccd1 vccd1 _2780_/D sky130_fd_sc_hd__and3_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1274_ _2193_/A vssd1 vssd1 vccd1 vccd1 _1299_/B sky130_fd_sc_hd__buf_1
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3013_ _3091_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3013_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_114_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2728_ _2728_/CLK _2728_/D vssd1 vssd1 vccd1 vccd1 _2728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput430 _2761_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__clkbuf_2
X_2659_ _1676_/Y _1709_/Y _1670_/Y _1728_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2659_/X sky130_fd_sc_hd__mux4_1
Xoutput441 _2737_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput452 _2356_/X vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput463 _2366_/X vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__clkbuf_2
Xoutput474 _2376_/X vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput485 _2237_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput496 _2247_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1961_ _2713_/Q _1961_/B vssd1 vssd1 vccd1 vccd1 _1962_/A sky130_fd_sc_hd__nand2_1
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1892_ _2692_/Q _1884_/X _2724_/Q _1887_/X vssd1 vssd1 vccd1 vccd1 _2692_/D sky130_fd_sc_hd__a22o_1
XFILLER_204_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2513_ _2512_/X _2778_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2444_ _2604_/X _2443_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2375_ _2754_/Q vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1326_ _2105_/A vssd1 vssd1 vccd1 vccd1 _1326_/X sky130_fd_sc_hd__buf_1
XFILLER_211_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1257_ _1285_/A _2203_/B _2642_/X vssd1 vssd1 vccd1 vccd1 _2768_/D sky130_fd_sc_hd__and3_1
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2160_ _3111_/Q _2147_/X _3033_/Q _2159_/X vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__a22o_1
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2091_ _2397_/S vssd1 vssd1 vccd1 vccd1 _2118_/B sky130_fd_sc_hd__inv_2
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2993_ _3110_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2993_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_72_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1944_ _1944_/A vssd1 vssd1 vccd1 vccd1 _1945_/B sky130_fd_sc_hd__inv_2
XFILLER_187_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1875_ _1878_/A _2456_/X vssd1 vssd1 vccd1 vccd1 _2701_/D sky130_fd_sc_hd__and2_1
XFILLER_175_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2427_ _2588_/X _2427_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2358_ _2737_/Q vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ _1319_/A _1333_/B _2649_/X vssd1 vssd1 vccd1 vccd1 _2775_/D sky130_fd_sc_hd__and3_1
XFILLER_211_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2289_ vssd1 vssd1 vccd1 vccd1 _2289_/HI _2289_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1660_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1665_/A sky130_fd_sc_hd__buf_1
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1591_ _1548_/B _1590_/X _1548_/B _1590_/X vssd1 vssd1 vccd1 vccd1 _1591_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2212_ vssd1 vssd1 vccd1 vccd1 _2212_/HI _2212_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2143_ _3070_/Q _2120_/X _2914_/Q _2124_/X vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2074_ _2081_/B vssd1 vssd1 vccd1 vccd1 _2080_/B sky130_fd_sc_hd__buf_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2976_ _3093_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2976_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_194_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1927_ _2667_/Q _1921_/X _2699_/Q _1922_/X vssd1 vssd1 vccd1 vccd1 _2667_/D sky130_fd_sc_hd__a22o_1
XFILLER_198_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1858_ _1860_/A _2420_/X vssd1 vssd1 vccd1 vccd1 _2715_/D sky130_fd_sc_hd__and2_1
XFILLER_190_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1789_ _2779_/Q _2777_/Q _1683_/Y _1727_/Y vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__o22a_1
XFILLER_150_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput330 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 _2447_/A1 sky130_fd_sc_hd__buf_1
XFILLER_27_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput341 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 _2449_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput352 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 _2451_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput363 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _2010_/B sky130_fd_sc_hd__clkbuf_1
XPHY_7384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2830_ _3103_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2830_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2761_ _2761_/CLK _2761_/D vssd1 vssd1 vccd1 vccd1 _2761_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1712_ _1707_/X _1711_/X _1707_/X _1711_/X vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2692_ _2729_/CLK _2692_/D vssd1 vssd1 vccd1 vccd1 _2692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_1 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _1647_/A _2522_/X vssd1 vssd1 vccd1 vccd1 _2749_/D sky130_fd_sc_hd__and2_1
XFILLER_103_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1574_ _1572_/Y _1573_/X _1572_/Y _1573_/X vssd1 vssd1 vccd1 vccd1 _1574_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2126_ _2950_/Q _2114_/X _2989_/Q _2117_/X _2125_/X vssd1 vssd1 vccd1 vccd1 _2126_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ _2065_/B _2078_/A vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__or2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2959_ _3076_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2959_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1290_ _2178_/A vssd1 vssd1 vccd1 vccd1 _1319_/A sky130_fd_sc_hd__buf_1
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput160 la_data_in[94] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_1
XFILLER_188_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput171 la_oenb[103] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__buf_1
XFILLER_49_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput182 la_oenb[113] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_hd__buf_1
Xinput193 la_oenb[123] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__buf_1
XFILLER_188_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2813_ _3086_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2813_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_73_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2744_ _2761_/CLK _2744_/D vssd1 vssd1 vccd1 vccd1 _2744_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2675_ _2722_/CLK _2675_/D vssd1 vssd1 vccd1 vccd1 _2675_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput601 _2668_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1626_ _1660_/A vssd1 vssd1 vccd1 vccd1 _2134_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_177_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1557_ _1445_/B _1465_/A _1527_/X _1466_/B vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1488_ _1490_/A _1488_/B vssd1 vssd1 vccd1 vccd1 _3102_/D sky130_fd_sc_hd__nor2_4
XFILLER_45_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2109_ _2109_/A vssd1 vssd1 vccd1 vccd1 _2109_/X sky130_fd_sc_hd__buf_1
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3089_ _3089_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3089_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2460_ _2619_/X _2459_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1411_ _2869_/Q _2102_/A _1408_/X _1410_/X vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__a211o_1
XFILLER_9_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2391_ _1400_/X _2828_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1342_ _2193_/A vssd1 vssd1 vccd1 vccd1 _1367_/B sky130_fd_sc_hd__buf_1
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1273_ _2848_/Q _1266_/X _1268_/X _1272_/X vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__a211o_1
XFILLER_211_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3012_ _3090_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3012_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2727_ _2729_/CLK _2727_/D vssd1 vssd1 vccd1 vccd1 _2727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput420 _2752_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2658_ _2655_/X _2656_/X _2657_/X _2626_/X _2053_/B _1834_/A vssd1 vssd1 vccd1 vccd1
+ _2658_/X sky130_fd_sc_hd__mux4_1
Xoutput431 _2209_/LO vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput442 _2738_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput453 _2357_/X vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput464 _2367_/X vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__clkbuf_2
X_1609_ _1607_/Y _1609_/B _1855_/A _1609_/D vssd1 vssd1 vccd1 vccd1 _3112_/D sky130_fd_sc_hd__and4b_4
X_2589_ _2008_/X _2720_/Q _2589_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__mux2_1
Xoutput475 _2377_/X vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__clkbuf_2
Xoutput486 _2219_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput497 _2220_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1960_ _1960_/A vssd1 vssd1 vccd1 vccd1 _1961_/B sky130_fd_sc_hd__inv_2
XFILLER_18_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1891_ _2693_/Q _1884_/X _2725_/Q _1887_/X vssd1 vssd1 vccd1 vccd1 _2693_/D sky130_fd_sc_hd__a22o_1
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2512_ _2511_/X _2778_/Q _2557_/S vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2443_ _2604_/X _2443_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2443_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2374_ _2753_/Q vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1325_ _1353_/A _1333_/B _2380_/X vssd1 vssd1 vccd1 vccd1 _2778_/D sky130_fd_sc_hd__and3_1
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1256_ _2178_/A vssd1 vssd1 vccd1 vccd1 _1285_/A sky130_fd_sc_hd__buf_1
XFILLER_84_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2090_ _2398_/S vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__inv_2
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2992_ _3109_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2992_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_128_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1943_ _2704_/Q _1943_/B vssd1 vssd1 vccd1 vccd1 _1944_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1874_ _1878_/A _2458_/X vssd1 vssd1 vccd1 vccd1 _2702_/D sky130_fd_sc_hd__and2_1
XFILLER_70_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2426_ _2586_/X _2425_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2357_ _2736_/Q vssd1 vssd1 vccd1 vccd1 _2357_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1308_ _2193_/A vssd1 vssd1 vccd1 vccd1 _1333_/B sky130_fd_sc_hd__buf_1
XFILLER_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2288_ vssd1 vssd1 vccd1 vccd1 _2288_/HI _2288_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1590_ _1569_/X _1589_/X _1569_/X _1589_/X vssd1 vssd1 vccd1 vccd1 _1590_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2211_ vssd1 vssd1 vccd1 vccd1 _2211_/HI _2211_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2142_ _3109_/Q _2106_/X _3031_/Q _2109_/X vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2073_ _2073_/A _2078_/B vssd1 vssd1 vccd1 vccd1 _2517_/S sky130_fd_sc_hd__or2_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2975_ _3092_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2975_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_194_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1926_ _2668_/Q _1921_/X _2700_/Q _1922_/X vssd1 vssd1 vccd1 vccd1 _2668_/D sky130_fd_sc_hd__a22o_1
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1857_ _1860_/A _2422_/X vssd1 vssd1 vccd1 vccd1 _2716_/D sky130_fd_sc_hd__and2_1
XFILLER_198_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1788_ _2798_/Q _1734_/Y _1787_/Y _2773_/Q vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__a22o_1
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2409_ _2570_/X _2409_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__mux2_1
XPHY_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput320 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 input320/X sky130_fd_sc_hd__buf_1
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput331 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 _2435_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_209_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput342 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 _2423_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput353 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 _2411_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput364 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _2001_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2760_ _2761_/CLK _2760_/D vssd1 vssd1 vccd1 vccd1 _2760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1711_ _2787_/Q _1708_/X _1709_/Y _1710_/Y vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__o22a_1
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2691_ _2722_/CLK _2691_/D vssd1 vssd1 vccd1 vccd1 _2691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_2 _2177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1642_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1647_/A sky130_fd_sc_hd__buf_1
XFILLER_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1573_ _1473_/B _1551_/A _1472_/A _1551_/Y vssd1 vssd1 vccd1 vccd1 _1573_/X sky130_fd_sc_hd__o22a_1
XFILLER_28_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2125_ _3067_/Q _2120_/X _2911_/Q _2124_/X vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2056_ _2060_/A _2079_/A vssd1 vssd1 vccd1 vccd1 _2487_/S sky130_fd_sc_hd__or2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2958_ _3075_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2958_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1909_ _2681_/Q _1907_/X _2713_/Q _1908_/X vssd1 vssd1 vccd1 vccd1 _2681_/D sky130_fd_sc_hd__a22o_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2889_ _3084_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2889_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_87_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput150 la_data_in[85] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__buf_1
XPHY_7171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput161 la_data_in[95] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_1
XFILLER_209_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput172 la_oenb[104] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_hd__buf_1
XPHY_7193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput183 la_oenb[114] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__buf_1
Xinput194 la_oenb[124] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__buf_1
XPHY_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2812_ _3085_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2812_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_158_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2743_ _2761_/CLK _2743_/D vssd1 vssd1 vccd1 vccd1 _2743_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_160_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2674_ _2722_/CLK _2674_/D vssd1 vssd1 vccd1 vccd1 _2674_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput602 _2669_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1625_ _2139_/A vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1556_ _1433_/B _1472_/A _1432_/A _1473_/B vssd1 vssd1 vccd1 vccd1 _1556_/X sky130_fd_sc_hd__o22a_1
XFILLER_138_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1487_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__inv_2
XFILLER_115_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2108_ _2158_/A vssd1 vssd1 vccd1 vccd1 _2109_/A sky130_fd_sc_hd__buf_1
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3088_ _3088_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3088_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2039_ _2047_/A _2088_/A vssd1 vssd1 vccd1 vccd1 _2466_/S sky130_fd_sc_hd__or2_1
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1410_ _2947_/Q _2114_/A _2986_/Q _2117_/A _1409_/X vssd1 vssd1 vccd1 vccd1 _1410_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2390_ _1391_/X _2827_/Q _2652_/S vssd1 vssd1 vccd1 vccd1 _2390_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1341_ _2858_/Q _1334_/X _1336_/X _1340_/X vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__a211o_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1272_ _2926_/Q _1269_/X _2965_/Q _1270_/X _1271_/X vssd1 vssd1 vccd1 vccd1 _1272_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _3089_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3011_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_209_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2726_ _2728_/CLK _2726_/D vssd1 vssd1 vccd1 vccd1 _2726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput410 _2743_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2657_ _1698_/Y _1673_/Y _1822_/Y _1684_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2657_/X sky130_fd_sc_hd__mux4_1
Xoutput421 _2753_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__clkbuf_2
Xoutput432 _2210_/LO vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput443 _2739_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1608_ _1608_/A _1608_/B vssd1 vssd1 vccd1 vccd1 _1609_/D sky130_fd_sc_hd__nand2_1
Xoutput454 _2358_/X vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__clkbuf_2
X_2588_ _2719_/Q _2587_/X _2621_/S vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
Xoutput465 _2368_/X vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput476 _2378_/X vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__clkbuf_2
Xoutput487 _2238_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput498 _2248_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1539_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1539_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1890_ _2694_/Q _1884_/X _2726_/Q _1887_/X vssd1 vssd1 vccd1 vccd1 _2694_/D sky130_fd_sc_hd__a22o_1
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2511_ _2628_/X _2778_/Q _2511_/S vssd1 vssd1 vccd1 vccd1 _2511_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2442_ _2602_/X _2441_/X _2462_/S vssd1 vssd1 vccd1 vccd1 _2442_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2373_ _2752_/Q vssd1 vssd1 vccd1 vccd1 _2373_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1324_ _2178_/A vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__buf_1
XFILLER_42_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1255_ _2846_/Q _2195_/X _1252_/X _1254_/X vssd1 vssd1 vccd1 vccd1 _1255_/X sky130_fd_sc_hd__a211o_1
XFILLER_204_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2709_ _2722_/CLK _2709_/D vssd1 vssd1 vccd1 vccd1 _2709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2991_ _3108_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2991_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1942_ _1942_/A vssd1 vssd1 vccd1 vccd1 _1943_/B sky130_fd_sc_hd__inv_2
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1873_ _2154_/A vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2425_ _2586_/X _2425_/A1 _2429_/S vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2356_ _2735_/Q vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1307_ _2853_/Q _1300_/X _1302_/X _1306_/X vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__a211o_1
XPHY_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2287_ vssd1 vssd1 vccd1 vccd1 _2287_/HI _2287_/LO sky130_fd_sc_hd__conb_1
XFILLER_38_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2210_ vssd1 vssd1 vccd1 vccd1 _2210_/HI _2210_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2141_ _2173_/A _2146_/B _2631_/X vssd1 vssd1 vccd1 vccd1 _2796_/D sky130_fd_sc_hd__and3_1
XFILLER_208_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2072_ _2072_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2514_/S sky130_fd_sc_hd__or2_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2974_ _3091_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2974_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_17_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1925_ _2669_/Q _1921_/X _2701_/Q _1922_/X vssd1 vssd1 vccd1 vccd1 _2669_/D sky130_fd_sc_hd__a22o_1
X_1856_ _1860_/A _2424_/X vssd1 vssd1 vccd1 vccd1 _2717_/D sky130_fd_sc_hd__and2_1
XFILLER_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1787_ _2798_/Q vssd1 vssd1 vccd1 vccd1 _1787_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2408_ _2568_/X _2407_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2339_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput310 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 input310/X sky130_fd_sc_hd__buf_1
XPHY_7331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput321 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 input321/X sky130_fd_sc_hd__buf_1
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput332 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 _2437_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput343 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 _2425_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_209_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput354 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 _2413_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput365 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1710_ _2791_/Q vssd1 vssd1 vccd1 vccd1 _1710_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2690_ _2722_/CLK _2690_/D vssd1 vssd1 vccd1 vccd1 _2690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1641_ _1641_/A _2525_/X vssd1 vssd1 vccd1 vccd1 _2750_/D sky130_fd_sc_hd__and2_1
XANTENNA_3 _2760_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1572_ _1572_/A vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2124_ _2188_/A vssd1 vssd1 vccd1 vccd1 _2124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2055_ _2061_/B _2078_/A vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__or2_1
XFILLER_208_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _3074_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2957_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1908_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1908_/X sky130_fd_sc_hd__buf_1
XFILLER_191_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2888_ _3083_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2888_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1839_ _2192_/A vssd1 vssd1 vccd1 vccd1 _2154_/A sky130_fd_sc_hd__buf_2
XFILLER_11_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput140 la_data_in[76] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__buf_1
XPHY_7161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput151 la_data_in[86] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__buf_1
XFILLER_49_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput162 la_data_in[96] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__buf_1
XPHY_7183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 la_oenb[105] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_hd__buf_1
XFILLER_209_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 la_oenb[115] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_hd__buf_1
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_oenb[125] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__buf_1
XFILLER_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2811_ _3084_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2811_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2742_ _2761_/CLK _2742_/D vssd1 vssd1 vccd1 vccd1 _2742_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _2722_/CLK _2673_/D vssd1 vssd1 vccd1 vccd1 _2673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput603 _2670_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_2
X_1624_ _2607_/S vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_126_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1555_ _1539_/Y _1554_/A _1539_/A _1554_/Y vssd1 vssd1 vccd1 vccd1 _1555_/X sky130_fd_sc_hd__o22a_1
XFILLER_154_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1486_ _1490_/A _1486_/B vssd1 vssd1 vccd1 vccd1 _3101_/D sky130_fd_sc_hd__nor2_4
XFILLER_119_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2107_ _2107_/A _2107_/B vssd1 vssd1 vccd1 vccd1 _2158_/A sky130_fd_sc_hd__nor2_2
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3087_ _3087_/D _1622_/X vssd1 vssd1 vccd1 vccd1 _3087_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2061_/B _2087_/A vssd1 vssd1 vccd1 vccd1 _2088_/A sky130_fd_sc_hd__or2_1
XFILLER_149_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ _2936_/Q _1337_/X _2975_/Q _1338_/X _1339_/X vssd1 vssd1 vccd1 vccd1 _1340_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1271_ _3043_/Q _1260_/X _2887_/Q _1261_/X vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3010_ _3088_/D _1620_/X vssd1 vssd1 vccd1 vccd1 _3010_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_37_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2725_ _2728_/CLK _2725_/D vssd1 vssd1 vccd1 vccd1 _2725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput400 _2319_/X vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__clkbuf_2
X_2656_ _1721_/Y _1666_/Y _1689_/Y _1678_/Y _2625_/S _2626_/S vssd1 vssd1 vccd1 vccd1
+ _2656_/X sky130_fd_sc_hd__mux4_1
Xoutput411 _2744_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput422 _2754_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput433 _2211_/LO vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1607_ _1608_/A _1608_/B vssd1 vssd1 vccd1 vccd1 _1607_/Y sky130_fd_sc_hd__nor2_1
Xoutput444 _2215_/LO vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__clkbuf_2
X_2587_ _2007_/X _2719_/Q _2620_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
Xoutput455 _2359_/X vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__clkbuf_2
Xoutput466 _2369_/X vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__clkbuf_2
Xoutput477 _2379_/X vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__clkbuf_2
X_1538_ _1441_/B _1537_/X _1441_/B _1537_/X vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__a2bb2o_2
Xoutput488 _2239_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput499 _2249_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1469_ _1480_/A vssd1 vssd1 vccd1 vccd1 _1479_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2510_ _2509_/X _2777_/Q _2558_/S vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2441_ _2602_/X _2441_/A1 _2445_/S vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2372_ _2751_/Q vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1323_ _2856_/Q _1300_/X _1320_/X _1322_/X vssd1 vssd1 vccd1 vccd1 _1323_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1254_ _2924_/Q _2198_/X _2963_/Q _2199_/X _1253_/X vssd1 vssd1 vccd1 vccd1 _1254_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2708_ _2722_/CLK _2708_/D vssd1 vssd1 vccd1 vccd1 _2708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2639_ _2202_/X _2804_/Q _2645_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2990_ _3107_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2990_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_91_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1941_ _2703_/Q _1941_/B vssd1 vssd1 vccd1 vccd1 _1942_/A sky130_fd_sc_hd__nand2_1
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1872_ _1872_/A _2460_/X vssd1 vssd1 vccd1 vccd1 _2703_/D sky130_fd_sc_hd__and2_1
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2424_ _2584_/X _2423_/X _2448_/S vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2355_ _2734_/Q vssd1 vssd1 vccd1 vccd1 _2355_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1306_ _2931_/Q _1303_/X _2970_/Q _1304_/X _1305_/X vssd1 vssd1 vccd1 vccd1 _1306_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2286_ vssd1 vssd1 vccd1 vccd1 _2286_/HI _2286_/LO sky130_fd_sc_hd__conb_1
XFILLER_168_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2140_ _2178_/A vssd1 vssd1 vccd1 vccd1 _2173_/A sky130_fd_sc_hd__buf_1
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2071_ _2089_/A _2072_/B vssd1 vssd1 vccd1 vccd1 _2511_/S sky130_fd_sc_hd__or2_1
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _3090_/D _1619_/X vssd1 vssd1 vccd1 vccd1 _2973_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1924_ _2670_/Q _1921_/X _2702_/Q _1922_/X vssd1 vssd1 vccd1 vccd1 _2670_/D sky130_fd_sc_hd__a22o_1
XFILLER_202_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1855_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1860_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1786_ _1706_/Y _2786_/Q _2782_/Q _1676_/Y vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2407_ _2568_/X _2407_/A1 _2413_/S vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2338_ _2350_/A vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2269_ vssd1 vssd1 vccd1 vccd1 _2269_/HI _2269_/LO sky130_fd_sc_hd__conb_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput300 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input300/X sky130_fd_sc_hd__buf_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput311 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 input311/X sky130_fd_sc_hd__buf_1
XFILLER_1_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput322 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input322/X sky130_fd_sc_hd__buf_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput333 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 _2439_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput344 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 _2427_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput355 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 _2453_/A1 sky130_fd_sc_hd__clkbuf_1
XPHY_7376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput366 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _1880_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1640_ _1641_/A _2528_/X vssd1 vssd1 vccd1 vccd1 _2751_/D sky130_fd_sc_hd__and2_1
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_4 _2761_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1571_ _1452_/B _1458_/A _1451_/A _1459_/B vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__o22a_1
XFILLER_67_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2123_ _2123_/A vssd1 vssd1 vccd1 vccd1 _2188_/A sky130_fd_sc_hd__buf_1
XFILLER_132_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2054_ _2087_/C _2054_/B _2078_/A vssd1 vssd1 vccd1 vccd1 _2484_/S sky130_fd_sc_hd__or3_1
XFILLER_78_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2956_ _3112_/D _1616_/X vssd1 vssd1 vccd1 vccd1 _2956_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_202_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1907_ _1921_/A vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2887_ _3082_/D _1615_/X vssd1 vssd1 vccd1 vccd1 _2887_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_191_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1838_ _1882_/A vssd1 vssd1 vccd1 vccd1 _2192_/A sky130_fd_sc_hd__buf_2
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1769_ _1767_/X _1768_/X _1767_/X _1768_/X vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput130 la_data_in[67] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__buf_1
XPHY_7151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput141 la_data_in[77] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_1
XFILLER_209_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput152 la_data_in[87] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_1
XPHY_7173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput163 la_data_in[97] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__buf_1
XPHY_7184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 la_oenb[106] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_hd__buf_1
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput185 la_oenb[116] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_1
XPHY_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 la_oenb[126] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__buf_1
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2810_ _3083_/D _1612_/Y vssd1 vssd1 vccd1 vccd1 _2810_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2741_ _2761_/CLK _2741_/D vssd1 vssd1 vccd1 vccd1 _2741_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_201_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2672_ _2722_/CLK _2672_/D vssd1 vssd1 vccd1 vccd1 _2672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1623_ _2134_/A _2558_/X vssd1 vssd1 vccd1 vccd1 _2761_/D sky130_fd_sc_hd__and2_2
Xoutput604 _2671_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1554_ _1554_/A vssd1 vssd1 vccd1 vccd1 _1554_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1485_ _1485_/A vssd1 vssd1 vccd1 vccd1 _1486_/B sky130_fd_sc_hd__inv_2
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

