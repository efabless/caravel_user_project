VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_32_256_sky130
   CLASS BLOCK ;
   SIZE 472.3 BY 219.34 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.88 0.0 113.26 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.32 0.0 118.7 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  124.44 0.0 124.82 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.88 0.0 130.26 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.0 0.0 136.38 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.8 0.0 143.18 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.56 0.0 147.94 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.12 0.0 159.5 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.24 0.0 165.62 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.8 0.0 177.18 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.92 0.0 183.3 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 0.0 195.54 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  200.6 0.0 200.98 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.72 0.0 207.1 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 0.0 213.22 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.08 0.0 242.46 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 0.0 247.9 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 0.0 253.34 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 0.0 259.46 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.2 0.0 265.58 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  270.64 0.0 271.02 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 0.0 282.58 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 0.0 288.02 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 0.0 294.82 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 0.0 299.58 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  77.52 0.0 77.9 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.64 0.0 84.02 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 132.6 0.38 132.98 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 140.76 0.38 141.14 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 146.88 0.38 147.26 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  67.32 218.96 67.7 219.34 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  66.64 218.96 67.02 219.34 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  65.96 218.96 66.34 219.34 ;
      END
   END addr0[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.72 0.38 37.1 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 45.56 0.38 45.94 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 37.4 0.38 37.78 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.76 0.0 90.14 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.2 0.0 95.58 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.0 0.0 102.38 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.44 0.0 107.82 0.38 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.0 0.0 306.38 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.92 0.0 149.3 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 0.0 189.42 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 0.0 198.94 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 0.0 216.62 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 0.0 239.06 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 0.0 268.98 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 0.0 289.38 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.92 0.0 319.3 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.12 0.0 329.5 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  338.64 0.0 339.02 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.84 0.0 349.22 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.04 0.0 359.42 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  369.24 0.0 369.62 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 0.0 377.78 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  388.96 0.0 389.34 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  399.16 0.0 399.54 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  408.68 0.0 409.06 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  471.92 58.48 472.3 58.86 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  471.92 59.16 472.3 59.54 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  471.92 63.92 472.3 64.3 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  471.92 59.84 472.3 60.22 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  471.92 61.88 472.3 62.26 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  469.2 1.36 470.94 217.98 ;
         LAYER met3 ;
         RECT  1.36 216.24 470.94 217.98 ;
         LAYER met3 ;
         RECT  1.36 1.36 470.94 3.1 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 217.98 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 214.58 ;
         LAYER met3 ;
         RECT  4.76 212.84 467.54 214.58 ;
         LAYER met3 ;
         RECT  4.76 4.76 467.54 6.5 ;
         LAYER met4 ;
         RECT  465.8 4.76 467.54 214.58 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 471.68 218.72 ;
   LAYER  met2 ;
      RECT  0.62 0.62 471.68 218.72 ;
   LAYER  met3 ;
      RECT  0.98 132.0 471.68 133.58 ;
      RECT  0.62 133.58 0.98 140.16 ;
      RECT  0.62 141.74 0.98 146.28 ;
      RECT  0.62 46.54 0.98 132.0 ;
      RECT  0.62 38.38 0.98 44.96 ;
      RECT  0.98 57.88 471.32 59.46 ;
      RECT  0.98 59.46 471.32 132.0 ;
      RECT  471.32 64.9 471.68 132.0 ;
      RECT  471.32 60.82 471.68 61.28 ;
      RECT  471.32 62.86 471.68 63.32 ;
      RECT  0.98 218.58 471.54 218.72 ;
      RECT  471.54 133.58 471.68 215.64 ;
      RECT  471.54 215.64 471.68 218.58 ;
      RECT  471.54 218.58 471.68 218.72 ;
      RECT  0.62 147.86 0.76 215.64 ;
      RECT  0.62 215.64 0.76 218.58 ;
      RECT  0.62 218.58 0.76 218.72 ;
      RECT  0.76 147.86 0.98 215.64 ;
      RECT  0.76 218.58 0.98 218.72 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 36.12 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 36.12 ;
      RECT  0.98 0.62 471.32 0.76 ;
      RECT  471.32 0.62 471.54 0.76 ;
      RECT  471.32 3.7 471.54 57.88 ;
      RECT  471.54 0.62 471.68 0.76 ;
      RECT  471.54 0.76 471.68 3.7 ;
      RECT  471.54 3.7 471.68 57.88 ;
      RECT  0.98 133.58 4.16 212.24 ;
      RECT  0.98 212.24 4.16 215.18 ;
      RECT  0.98 215.18 4.16 215.64 ;
      RECT  4.16 133.58 468.14 212.24 ;
      RECT  4.16 215.18 468.14 215.64 ;
      RECT  468.14 133.58 471.54 212.24 ;
      RECT  468.14 212.24 471.54 215.18 ;
      RECT  468.14 215.18 471.54 215.64 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 57.88 ;
      RECT  4.16 3.7 468.14 4.16 ;
      RECT  4.16 7.1 468.14 57.88 ;
      RECT  468.14 3.7 471.32 4.16 ;
      RECT  468.14 4.16 471.32 7.1 ;
      RECT  468.14 7.1 471.32 57.88 ;
   LAYER  met4 ;
      RECT  112.28 0.98 113.86 218.72 ;
      RECT  113.86 0.62 117.72 0.98 ;
      RECT  119.3 0.62 123.84 0.98 ;
      RECT  125.42 0.62 129.28 0.98 ;
      RECT  130.86 0.62 135.4 0.98 ;
      RECT  143.78 0.62 146.96 0.98 ;
      RECT  160.1 0.62 164.64 0.98 ;
      RECT  171.66 0.62 176.2 0.98 ;
      RECT  183.9 0.62 187.76 0.98 ;
      RECT  201.58 0.62 206.12 0.98 ;
      RECT  218.58 0.62 223.8 0.98 ;
      RECT  230.82 0.62 235.36 0.98 ;
      RECT  243.06 0.62 246.92 0.98 ;
      RECT  260.06 0.62 264.6 0.98 ;
      RECT  271.62 0.62 275.48 0.98 ;
      RECT  283.18 0.62 287.04 0.98 ;
      RECT  78.5 0.62 83.04 0.98 ;
      RECT  66.72 0.98 68.3 218.36 ;
      RECT  68.3 0.98 112.28 218.36 ;
      RECT  68.3 218.36 112.28 218.72 ;
      RECT  84.62 0.62 89.16 0.98 ;
      RECT  90.74 0.62 94.6 0.98 ;
      RECT  96.18 0.62 101.4 0.98 ;
      RECT  102.98 0.62 106.84 0.98 ;
      RECT  108.42 0.62 112.28 0.98 ;
      RECT  300.18 0.62 305.4 0.98 ;
      RECT  136.98 0.62 138.8 0.98 ;
      RECT  140.38 0.62 142.2 0.98 ;
      RECT  149.9 0.62 153.08 0.98 ;
      RECT  154.66 0.62 157.16 0.98 ;
      RECT  166.22 0.62 168.04 0.98 ;
      RECT  169.62 0.62 170.08 0.98 ;
      RECT  177.78 0.62 178.24 0.98 ;
      RECT  179.82 0.62 182.32 0.98 ;
      RECT  190.02 0.62 194.56 0.98 ;
      RECT  196.14 0.62 197.96 0.98 ;
      RECT  199.54 0.62 200.0 0.98 ;
      RECT  207.7 0.62 208.16 0.98 ;
      RECT  209.74 0.62 212.24 0.98 ;
      RECT  213.82 0.62 215.64 0.98 ;
      RECT  225.38 0.62 227.2 0.98 ;
      RECT  228.78 0.62 229.24 0.98 ;
      RECT  236.94 0.62 238.08 0.98 ;
      RECT  239.66 0.62 241.48 0.98 ;
      RECT  249.86 0.62 252.36 0.98 ;
      RECT  253.94 0.62 256.44 0.98 ;
      RECT  258.02 0.62 258.48 0.98 ;
      RECT  266.18 0.62 268.0 0.98 ;
      RECT  269.58 0.62 270.04 0.98 ;
      RECT  277.06 0.62 278.2 0.98 ;
      RECT  279.78 0.62 281.6 0.98 ;
      RECT  289.98 0.62 293.84 0.98 ;
      RECT  295.42 0.62 297.24 0.98 ;
      RECT  306.98 0.62 308.8 0.98 ;
      RECT  310.38 0.62 318.32 0.98 ;
      RECT  319.9 0.62 328.52 0.98 ;
      RECT  330.1 0.62 338.04 0.98 ;
      RECT  339.62 0.62 348.24 0.98 ;
      RECT  349.82 0.62 358.44 0.98 ;
      RECT  360.02 0.62 368.64 0.98 ;
      RECT  370.22 0.62 376.8 0.98 ;
      RECT  378.38 0.62 388.36 0.98 ;
      RECT  389.94 0.62 398.56 0.98 ;
      RECT  400.14 0.62 408.08 0.98 ;
      RECT  113.86 218.58 468.6 218.72 ;
      RECT  468.6 218.58 471.54 218.72 ;
      RECT  471.54 0.98 471.68 218.58 ;
      RECT  471.54 218.58 471.68 218.72 ;
      RECT  409.66 0.62 468.6 0.76 ;
      RECT  409.66 0.76 468.6 0.98 ;
      RECT  468.6 0.62 471.54 0.76 ;
      RECT  471.54 0.62 471.68 0.76 ;
      RECT  471.54 0.76 471.68 0.98 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 76.92 0.76 ;
      RECT  3.7 0.76 76.92 0.98 ;
      RECT  0.62 0.98 0.76 218.36 ;
      RECT  0.62 218.36 0.76 218.58 ;
      RECT  0.62 218.58 0.76 218.72 ;
      RECT  0.76 218.58 3.7 218.72 ;
      RECT  3.7 218.36 65.36 218.58 ;
      RECT  3.7 218.58 65.36 218.72 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 215.18 ;
      RECT  3.7 215.18 4.16 218.36 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 215.18 7.1 218.36 ;
      RECT  7.1 0.98 66.72 4.16 ;
      RECT  7.1 4.16 66.72 215.18 ;
      RECT  7.1 215.18 66.72 218.36 ;
      RECT  113.86 0.98 465.2 4.16 ;
      RECT  113.86 4.16 465.2 215.18 ;
      RECT  113.86 215.18 465.2 218.58 ;
      RECT  465.2 0.98 468.14 4.16 ;
      RECT  465.2 215.18 468.14 218.58 ;
      RECT  468.14 0.98 468.6 4.16 ;
      RECT  468.14 4.16 468.6 215.18 ;
      RECT  468.14 215.18 468.6 218.58 ;
   END
END    sram_1rw0r0w_32_256_sky130
END    LIBRARY
