* SPICE3 file created from sparse_decoder.ext - technology: sky130A

.option scale=10000u

X0 m1_1250_153# li_23_n3860# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X1 decoder_cell_0_0[0]/a_12_n1# li_23_n3860# decoder_cell_0_0[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X2 m1_1250_153# li_235_204# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X3 decoder_cell_0_0[1]/a_12_n1# li_235_204# decoder_cell_0_0[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X4 m1_1250_153# li_448_n3912# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X5 decoder_cell_0_0[2]/a_12_n1# li_448_n3912# decoder_cell_0_0[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X6 m1_1250_153# li_659_202# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X7 decoder_cell_0_3[0]/a_12_n1# li_659_202# decoder_cell_0_0[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X8 m1_1233_n96# li_23_n3860# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X9 decoder_cell_0_1[0]/a_12_n1# li_23_n3860# decoder_cell_0_1[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X10 m1_1233_n96# li_235_204# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X11 decoder_cell_0_1[1]/a_12_n1# li_235_204# decoder_cell_0_1[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X12 m1_1233_n96# li_448_n3912# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X13 decoder_cell_0_1[2]/a_12_n1# li_448_n3912# decoder_cell_0_1[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X14 m1_1233_n96# li_659_202# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X15 decoder_cell_0_4/a_12_n1# li_659_202# decoder_cell_0_1[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X16 a_1331_n361# li_23_n3860# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X17 decoder_cell_0_2[0]/a_12_n1# li_23_n3860# decoder_cell_0_2[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X18 a_1331_n361# li_235_204# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X19 decoder_cell_0_2[1]/a_12_n1# li_235_204# decoder_cell_0_2[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X20 a_1331_n361# li_448_n3912# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X21 decoder_cell_0_6[0]/a_12_n1# li_448_n3912# decoder_cell_0_2[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X22 m1_1250_153# li_981_n3852# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X23 decoder_cell_0_3[0]/a_12_n1# li_981_n3852# decoder_cell_0_3[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X24 m1_1250_153# li_1189_223# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X25 decoder_cell_0_3[1]/a_12_n1# li_1189_223# m1_1250_153# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X26 m1_1233_n96# li_981_n3852# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X27 decoder_cell_0_4/a_12_n1# li_981_n3852# decoder_cell_0_5/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X28 m1_1233_n96# li_1081_202# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X29 m1_1233_n96# li_1081_202# decoder_cell_0_5/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X30 a_1331_n361# li_761_202# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X31 decoder_cell_0_6[0]/a_12_n1# li_761_202# decoder_cell_0_6[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X32 a_1331_n361# li_981_n3852# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X33 decoder_cell_0_6[1]/a_12_n1# li_981_n3852# decoder_cell_0_7/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X34 a_1331_n361# li_1081_202# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X35 a_1331_n361# li_1081_202# decoder_cell_0_7/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X36 a_1331_n459# li_23_n3860# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X37 decoder_cell_0_8[0]/a_12_n1# li_23_n3860# decoder_cell_0_8[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X38 a_1331_n459# li_235_204# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X39 decoder_cell_0_9[0]/a_12_n1# li_235_204# decoder_cell_0_8[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X40 a_1331_n459# li_549_n3836# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X41 decoder_cell_0_9[0]/a_12_n1# li_549_n3836# decoder_cell_0_9[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X42 a_1331_n459# li_761_202# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X43 decoder_cell_0_9[1]/a_12_n1# li_761_202# decoder_cell_0_10/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X44 a_1331_n3259# li_131_n3837# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X45 decoder_cell_0_60/a_12_n1# li_131_n3837# decoder_cell_0_60/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X46 a_1331_n2859# li_235_204# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X47 decoder_cell_0_50/a_12_n1# li_235_204# decoder_cell_0_50/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X48 a_1331_n3259# li_235_204# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X49 decoder_cell_0_61[0]/a_12_n1# li_235_204# decoder_cell_0_60/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X50 a_1331_n3259# li_448_n3912# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X51 decoder_cell_0_61[1]/a_12_n1# li_448_n3912# decoder_cell_0_61[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X52 li_23_n3860# buffer_0/li_48_5# buffer_0/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X53 li_23_n3860# buffer_0/li_48_5# buffer_0/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X54 li_131_n3837# li_23_n3860# buffer_0/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X55 li_131_n3837# li_23_n3860# buffer_0/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X56 a_1331_n2459# li_659_202# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X57 decoder_cell_0_40[0]/a_12_n1# li_659_202# decoder_cell_0_40[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X58 a_1331_n2459# li_869_n3865# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X59 decoder_cell_0_41/a_12_n1# li_869_n3865# decoder_cell_0_40[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X60 a_1331_n3161# li_869_n3865# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X61 decoder_cell_0_52/a_12_n1# li_869_n3865# decoder_cell_0_51/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X62 a_1331_n3561# li_659_202# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X63 decoder_cell_0_62/a_12_n1# li_659_202# decoder_cell_0_62/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X64 li_869_n3865# buffer_2/li_48_5# buffer_2/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X65 li_869_n3865# buffer_2/li_48_5# buffer_2/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X66 li_981_n3852# li_869_n3865# buffer_2/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X67 li_981_n3852# li_869_n3865# buffer_2/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X68 li_448_n3912# buffer_1/li_48_5# buffer_1/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X69 li_448_n3912# buffer_1/li_48_5# buffer_1/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X70 li_549_n3836# li_448_n3912# buffer_1/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X71 li_549_n3836# li_448_n3912# buffer_1/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X72 li_235_204# buffer_3/li_48_5# buffer_3/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X73 li_235_204# buffer_3/li_48_5# buffer_3/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X74 li_337_196# li_235_204# buffer_3/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X75 li_337_196# li_235_204# buffer_3/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X76 a_1329_n1961# li_448_n3912# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X77 decoder_cell_0_30[0]/a_12_n1# li_448_n3912# decoder_cell_0_33/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X78 a_1329_n1961# li_659_202# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X79 decoder_cell_0_30[1]/a_12_n1# li_659_202# decoder_cell_0_30[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X80 a_1329_n1961# li_869_n3865# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X81 decoder_cell_0_30[2]/a_12_n1# li_869_n3865# decoder_cell_0_30[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X82 a_1329_n1961# li_1081_202# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X83 a_1329_n1961# li_1081_202# decoder_cell_0_30[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X84 a_1331_n2459# li_1189_223# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X85 decoder_cell_0_41/a_12_n1# li_1189_223# a_1331_n2459# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X86 a_1331_n3161# li_1189_223# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X87 decoder_cell_0_52/a_12_n1# li_1189_223# a_1331_n3161# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X88 a_1331_n3659# li_659_202# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X89 decoder_cell_0_63/a_12_n1# li_659_202# decoder_cell_0_63/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X90 li_659_202# buffer_4/li_48_5# buffer_4/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X91 li_659_202# buffer_4/li_48_5# buffer_4/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X92 li_761_202# li_659_202# buffer_4/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X93 li_761_202# li_659_202# buffer_4/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X94 a_1331_n459# li_869_n3865# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X95 decoder_cell_0_11/a_12_n1# li_869_n3865# decoder_cell_0_10/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X96 a_1330_n1161# li_1189_223# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X97 decoder_cell_0_21/a_12_n1# li_1189_223# a_1330_n1161# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X98 a_1330_n1161# li_659_202# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X99 decoder_cell_0_20[0]/a_12_n1# li_659_202# decoder_cell_0_20[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X100 a_1330_n1161# li_869_n3865# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X101 decoder_cell_0_21/a_12_n1# li_869_n3865# decoder_cell_0_20[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X102 a_1329_n1961# li_131_n3837# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X103 decoder_cell_0_31/a_12_n1# li_131_n3837# decoder_cell_0_33/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X104 a_1329_n2059# li_131_n3837# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X105 decoder_cell_0_32/a_12_n1# li_131_n3837# decoder_cell_0_32/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X106 a_1331_n2761# li_549_n3836# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X107 decoder_cell_0_44/a_12_n1# li_549_n3836# decoder_cell_0_47/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X108 a_1331_n2859# li_549_n3836# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X109 decoder_cell_0_50/a_12_n1# li_549_n3836# decoder_cell_0_43[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X110 a_1331_n2859# li_761_202# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X111 decoder_cell_0_43[1]/a_12_n1# li_761_202# decoder_cell_0_43[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X112 a_1331_n2859# li_981_n3852# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X113 decoder_cell_0_43[2]/a_12_n1# li_981_n3852# decoder_cell_0_43[3]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X114 a_1331_n2859# li_1189_223# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X115 decoder_cell_0_43[3]/a_12_n1# li_1189_223# a_1331_n2859# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X116 a_1331_n3259# li_1081_202# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X117 a_1331_n3259# li_1081_202# decoder_cell_0_54/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X118 a_1331_n3259# li_761_202# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X119 decoder_cell_0_61[1]/a_12_n1# li_761_202# decoder_cell_0_53[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X120 a_1331_n3259# li_981_n3852# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X121 decoder_cell_0_53[1]/a_12_n1# li_981_n3852# decoder_cell_0_54/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X122 a_1331_n3659# li_131_n3837# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X123 decoder_cell_0_64/a_12_n1# li_131_n3837# decoder_cell_0_64/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X124 a_1331_n3659# li_235_204# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X125 decoder_cell_0_65[0]/a_12_n1# li_235_204# decoder_cell_0_64/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X126 a_1331_n3659# li_448_n3912# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X127 decoder_cell_0_63/a_n31_n1# li_448_n3912# decoder_cell_0_65[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X128 li_1081_202# buffer_5/li_48_5# buffer_5/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X129 li_1081_202# buffer_5/li_48_5# buffer_5/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X130 li_1189_223# li_1081_202# buffer_5/a_183_44# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X131 li_1189_223# li_1081_202# buffer_5/a_183_139# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X132 a_1331_n459# li_1189_223# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X133 decoder_cell_0_11/a_12_n1# li_1189_223# a_1331_n459# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X134 a_1330_n1259# li_23_n3860# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X135 decoder_cell_0_22/a_12_n1# li_23_n3860# decoder_cell_0_22/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X136 a_1329_n1961# li_337_196# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X137 decoder_cell_0_33/a_12_n1# li_337_196# decoder_cell_0_33/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X138 a_1331_n2761# li_235_204# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X139 decoder_cell_0_44/a_12_n1# li_235_204# decoder_cell_0_45/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X140 a_1331_n3161# li_131_n3837# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X141 decoder_cell_0_55/a_12_n1# li_131_n3837# decoder_cell_0_56/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X142 a_1331_n3561# li_235_204# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X143 decoder_cell_0_66[0]/a_12_n1# li_235_204# decoder_cell_0_67/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X144 a_1331_n3561# li_448_n3912# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X145 decoder_cell_0_62/a_n31_n1# li_448_n3912# decoder_cell_0_66[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X146 inv_lp_0/a_4_2# m1_1250_153# inv_lp_1/a_n39_2# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X147 inv_lp_0/a_4_2# m1_1250_153# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X148 a_1331_n761# li_23_n3860# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X149 decoder_cell_0_12[0]/a_12_n1# li_23_n3860# decoder_cell_0_12[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X150 a_1331_n761# li_235_204# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X151 decoder_cell_0_13[0]/a_12_n1# li_235_204# decoder_cell_0_12[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X152 a_1330_n1259# li_337_196# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X153 decoder_cell_0_22/a_12_n1# li_337_196# decoder_cell_0_23[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X154 a_1330_n1259# li_549_n3836# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X155 decoder_cell_0_23[1]/a_12_n1# li_549_n3836# decoder_cell_0_23[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X156 a_1330_n1259# li_761_202# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X157 decoder_cell_0_23[2]/a_12_n1# li_761_202# decoder_cell_0_23[3]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X158 a_1330_n1259# li_981_n3852# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X159 decoder_cell_0_23[3]/a_12_n1# li_981_n3852# decoder_cell_0_23[4]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X160 a_1330_n1259# li_1189_223# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X161 decoder_cell_0_23[4]/a_12_n1# li_1189_223# a_1330_n1259# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X162 a_1329_n2059# li_337_196# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X163 decoder_cell_0_32/a_n31_n1# li_337_196# decoder_cell_0_34[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X164 a_1329_n2059# li_549_n3836# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X165 decoder_cell_0_34[1]/a_12_n1# li_549_n3836# decoder_cell_0_34[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X166 a_1329_n2059# li_761_202# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X167 decoder_cell_0_34[2]/a_12_n1# li_761_202# decoder_cell_0_35[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X168 a_1331_n2761# li_131_n3837# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X169 decoder_cell_0_45/a_12_n1# li_131_n3837# decoder_cell_0_45/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X170 a_1331_n3161# li_235_204# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X171 decoder_cell_0_56/a_12_n1# li_235_204# decoder_cell_0_56/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X172 a_1331_n3561# li_131_n3837# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X173 decoder_cell_0_67/a_12_n1# li_131_n3837# decoder_cell_0_67/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X174 inv_lp_1/a_4_2# m1_1233_n96# inv_lp_1/a_n39_2# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X175 inv_lp_1/a_4_2# m1_1233_n96# m1_1269_0# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X176 a_1331_n761# li_549_n3836# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X177 decoder_cell_0_13[0]/a_12_n1# li_549_n3836# decoder_cell_0_13[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X178 a_1331_n761# li_761_202# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X179 decoder_cell_0_13[1]/a_12_n1# li_761_202# decoder_cell_0_13[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X180 a_1331_n761# li_981_n3852# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X181 decoder_cell_0_13[2]/a_12_n1# li_981_n3852# decoder_cell_0_13[3]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X182 a_1331_n761# li_1189_223# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X183 decoder_cell_0_13[3]/a_12_n1# li_1189_223# a_1331_n761# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X184 a_1331_n1561# li_23_n3860# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X185 decoder_cell_0_24/a_12_n1# li_23_n3860# decoder_cell_0_24/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X186 a_1329_n2059# li_869_n3865# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X187 decoder_cell_0_35[0]/a_12_n1# li_869_n3865# decoder_cell_0_35[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X188 a_1329_n2059# li_1081_202# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X189 a_1329_n2059# li_1081_202# decoder_cell_0_35[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X190 a_1331_n2761# li_981_n3852# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X191 decoder_cell_0_47/a_12_n1# li_981_n3852# decoder_cell_0_46[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X192 a_1331_n2761# li_1189_223# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X193 decoder_cell_0_46[1]/a_12_n1# li_1189_223# a_1331_n2761# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X194 a_1331_n3561# li_981_n3852# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X195 decoder_cell_0_62/a_12_n1# li_981_n3852# decoder_cell_0_58/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X196 a_1331_n859# li_23_n3860# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X197 decoder_cell_0_14[0]/a_12_n1# li_23_n3860# decoder_cell_0_14[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X198 a_1331_n859# li_235_204# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X199 decoder_cell_0_15/a_12_n1# li_235_204# decoder_cell_0_14[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X200 a_1331_n1561# li_337_196# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X201 decoder_cell_0_24/a_12_n1# li_337_196# decoder_cell_0_25[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X202 a_1331_n1561# li_549_n3836# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X203 decoder_cell_0_25[1]/a_12_n1# li_549_n3836# decoder_cell_0_25[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X204 a_1331_n1561# li_761_202# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X205 decoder_cell_0_25[2]/a_12_n1# li_761_202# decoder_cell_0_26[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X206 a_1331_n2361# li_337_196# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X207 decoder_cell_0_37/a_n31_n1# li_337_196# decoder_cell_0_36[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X208 a_1331_n2361# li_549_n3836# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X209 decoder_cell_0_36[1]/a_12_n1# li_549_n3836# decoder_cell_0_36[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X210 a_1331_n2361# li_761_202# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X211 decoder_cell_0_36[2]/a_12_n1# li_761_202# decoder_cell_0_36[3]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X212 a_1331_n2361# li_981_n3852# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X213 decoder_cell_0_36[3]/a_12_n1# li_981_n3852# decoder_cell_0_36[4]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X214 a_1331_n2361# li_1189_223# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X215 decoder_cell_0_36[4]/a_12_n1# li_1189_223# a_1331_n2361# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X216 a_1331_n2761# li_659_202# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X217 decoder_cell_0_47/a_12_n1# li_659_202# decoder_cell_0_47/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X218 a_1331_n3561# li_1081_202# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X219 a_1331_n3561# li_1081_202# decoder_cell_0_58/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X220 a_1331_n859# li_549_n3836# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X221 decoder_cell_0_15/a_12_n1# li_549_n3836# decoder_cell_0_16/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X222 a_1331_n1561# li_869_n3865# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X223 decoder_cell_0_26[0]/a_12_n1# li_869_n3865# decoder_cell_0_26[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X224 a_1331_n1561# li_1081_202# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X225 a_1331_n1561# li_1081_202# decoder_cell_0_26[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X226 a_1331_n2361# li_131_n3837# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X227 decoder_cell_0_37/a_12_n1# li_131_n3837# decoder_cell_0_37/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X228 a_1331_n3161# li_549_n3836# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X229 decoder_cell_0_56/a_12_n1# li_549_n3836# decoder_cell_0_48[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X230 a_1331_n3161# li_761_202# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X231 decoder_cell_0_48[1]/a_12_n1# li_761_202# decoder_cell_0_51/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X232 a_1331_n3659# li_981_n3852# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X233 decoder_cell_0_63/a_12_n1# li_981_n3852# decoder_cell_0_59[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X234 a_1331_n3659# li_1189_223# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X235 decoder_cell_0_59[1]/a_12_n1# li_1189_223# a_1331_n3659# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X236 a_1331_n859# li_659_202# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X237 decoder_cell_0_16/a_12_n1# li_659_202# decoder_cell_0_16/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X238 a_1331_n1659# li_23_n3860# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X239 decoder_cell_0_28/a_12_n1# li_23_n3860# decoder_cell_0_27/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X240 a_1331_n2459# li_131_n3837# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X241 decoder_cell_0_38/a_12_n1# li_131_n3837# decoder_cell_0_38/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X242 a_1331_n2859# li_131_n3837# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X243 decoder_cell_0_49/a_12_n1# li_131_n3837# decoder_cell_0_50/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X244 a_1331_n859# li_981_n3852# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X245 decoder_cell_0_16/a_12_n1# li_981_n3852# decoder_cell_0_17[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X246 a_1331_n859# li_1189_223# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X247 decoder_cell_0_17[1]/a_12_n1# li_1189_223# a_1331_n859# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X248 a_1330_n1161# li_23_n3860# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X249 decoder_cell_0_18/a_12_n1# li_23_n3860# decoder_cell_0_18/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X250 a_1331_n1659# li_448_n3912# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X251 decoder_cell_0_29[0]/a_12_n1# li_448_n3912# decoder_cell_0_28/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X252 a_1331_n1659# li_659_202# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X253 decoder_cell_0_29[1]/a_12_n1# li_659_202# decoder_cell_0_29[0]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X254 a_1331_n1659# li_869_n3865# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X255 decoder_cell_0_29[2]/a_12_n1# li_869_n3865# decoder_cell_0_29[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X256 a_1331_n1659# li_1081_202# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X257 a_1331_n1659# li_1081_202# decoder_cell_0_29[2]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X258 a_1331_n1659# li_337_196# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X259 decoder_cell_0_28/a_12_n1# li_337_196# decoder_cell_0_28/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X260 a_1331_n2459# li_337_196# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X261 decoder_cell_0_38/a_n31_n1# li_337_196# decoder_cell_0_39[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X262 a_1331_n2459# li_549_n3836# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X263 decoder_cell_0_39[1]/a_12_n1# li_549_n3836# decoder_cell_0_40[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X264 a_1330_n1161# li_337_196# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X265 decoder_cell_0_18/a_12_n1# li_337_196# decoder_cell_0_19[1]/a_12_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X266 a_1330_n1161# li_549_n3836# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X267 decoder_cell_0_19[1]/a_12_n1# li_549_n3836# decoder_cell_0_20[0]/a_n31_n1# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X268 a_1382_n334# a_1331_n361# a_1382_n432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X269 a_1382_n432# a_1331_n459# a_1382_n475# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X270 a_1382_n3534# a_1331_n3561# a_1477_n3632# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X271 a_1477_n3632# a_1331_n3659# a_1382_n3675# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X272 a_1382_n1534# a_1331_n1561# a_1477_n1632# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X273 a_1477_n1632# a_1331_n1659# a_1382_n1675# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X274 a_1382_n3534# a_1331_n3561# a_1382_n3632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X275 a_1382_n3632# a_1331_n3659# a_1382_n3675# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X276 a_1382_n1534# a_1331_n1561# a_1382_n1632# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X277 a_1382_n1632# a_1331_n1659# a_1382_n1675# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X278 a_1382_n3134# a_1331_n3161# a_1477_n3232# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X279 a_1477_n3232# a_1331_n3259# a_1382_n3275# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X280 a_1382_n3134# a_1331_n3161# a_1382_n3232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X281 a_1382_n3232# a_1331_n3259# a_1382_n3275# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X282 a_1382_n2734# a_1331_n2761# a_1477_n2832# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X283 a_1477_n2832# a_1331_n2859# a_1382_n2875# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X284 a_1380_n1934# a_1329_n1961# a_1475_n2032# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X285 a_1475_n2032# a_1329_n2059# a_1380_n2075# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X286 a_1380_n1934# a_1329_n1961# a_1380_n2032# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X287 a_1382_n2734# a_1331_n2761# a_1382_n2832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X288 a_1382_n2832# a_1331_n2859# a_1382_n2875# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X289 a_1381_n1134# a_1330_n1161# a_1476_n1232# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X290 a_1476_n1232# a_1330_n1259# a_1381_n1275# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X291 a_1380_n2032# a_1329_n2059# a_1380_n2075# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X292 a_1382_n2334# a_1331_n2361# a_1477_n2432# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X293 a_1477_n2432# a_1331_n2459# a_1382_n2475# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X294 a_1382_n734# a_1331_n761# a_1477_n832# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X295 a_1382_n734# a_1331_n761# a_1382_n832# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X296 a_1477_n832# a_1331_n859# a_1382_n875# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X297 a_1382_n832# a_1331_n859# a_1382_n875# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X298 a_1381_n1134# a_1330_n1161# a_1381_n1232# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X299 a_1381_n1232# a_1330_n1259# a_1381_n1275# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X300 a_1382_n2334# a_1331_n2361# a_1382_n2432# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X301 a_1382_n2432# a_1331_n2459# a_1382_n2475# w_1253_5# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X302 a_1382_n334# a_1331_n361# a_1477_n432# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
X303 a_1477_n432# a_1331_n459# a_1382_n475# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=15
C0 a_1382_n1632# SUB 3.00fF
C1 li_1189_223# SUB 6.76fF
C2 li_1081_202# SUB 7.57fF
C3 a_1382_n832# SUB 2.07fF
C4 li_337_196# SUB 6.83fF
C5 li_235_204# SUB 7.93fF
C6 a_1382_n3632# SUB 2.79fF
C7 a_1382_n3232# SUB 2.96fF
C8 a_1382_n2832# SUB 2.75fF
C9 a_1380_n2032# SUB 2.18fF
C10 li_549_n3836# SUB 7.08fF
C11 li_448_n3912# SUB 7.60fF
C12 li_981_n3852# SUB 7.14fF
C13 li_869_n3865# SUB 7.56fF
C14 li_761_202# SUB 6.99fF
C15 li_659_202# SUB 7.76fF
C16 a_1382_n2432# SUB 2.94fF
C17 li_131_n3837# SUB 6.96fF
C18 li_23_n3860# SUB 7.72fF
C19 w_1253_5# SUB 34.80fF
C20 a_1331_n459# SUB 2.01fF
C21 a_1382_n432# SUB 2.96fF
C22 a_1331_n361# SUB 2.02fF
C23 m1_1269_0# SUB 3.04fF
