`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***

//***Module***
module state_counters #(
        parameter integer WORD_SIZE = 32
    )
    (
        input  clk_i ,
        input  rst_i ,
        input  valid_i, 
        input  [3 : 0] wstrb_i,
        input  [WORD_SIZE -1 : 0] wdata_i,
        input  [1 : 0] operation_result_i ,
        input  valid_output_i,
        output  ready_o,
        output [WORD_SIZE - 1 : 0] rdata_o
    );

//***Internal logic generated by compiler***  


//***Dumped Internal logic***
    reg [WORD_SIZE-1:0] ecc_corrected_errors;
    reg [WORD_SIZE-1:0] ecc_uncorrected_errors;
    reg [WORD_SIZE-1:0] total_reads;
    reg ready_o;
    reg [WORD_SIZE-1:0] rdata_o;


    always @(posedge clk_i) begin

        if(rst_i) begin
            total_reads <= {WORD_SIZE {1'b0}}; 
            ecc_uncorrected_errors <= {WORD_SIZE {1'b0}}; 
            ecc_corrected_errors <= {WORD_SIZE {1'b0}}; 
        end
        else begin
            if (valid_output_i == 1'b1) begin
                total_reads <= total_reads +1;
                if (operation_result_i[0] == 1'b1) begin
                    ecc_corrected_errors <= ecc_corrected_errors + 1;
                end
                if (operation_result_i[1] == 1'b1) begin
                    ecc_uncorrected_errors <= ecc_uncorrected_errors + 1;
                end
            end
            if (valid_i) begin
                ready_o <= 1'b1;
                rdata_o = ecc_corrected_errors;
                if (wstrb_i[0]) ecc_corrected_errors[7:0]   <= wdata_i[7:0];
                if (wstrb_i[1]) ecc_corrected_errors[15:8]  <= wdata_i[15:8];
                if (wstrb_i[2]) ecc_corrected_errors[23:16] <= wdata_i[23:16];
                if (wstrb_i[3]) ecc_corrected_errors[31:24] <= wdata_i[31:24];
            end
        end
    end

    
//***Handcrafted Internal logic*** 
//TODO
endmodule
