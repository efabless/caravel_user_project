magic
tech sky130A
magscale 1 2
timestamp 1640845691
<< nwell >>
rect -186 182 976 358
<< nmos >>
rect -10 -124 26 -40
rect 84 -124 120 -40
rect 214 -124 250 -40
rect 352 -124 388 -40
rect 446 -124 482 -40
rect 648 -124 684 -40
rect 746 -124 782 -40
<< pmos >>
rect -10 226 26 310
rect 84 226 120 310
rect 214 226 250 310
rect 352 226 388 310
rect 658 226 694 310
rect 752 226 788 310
<< ndiff >>
rect -64 -64 -10 -40
rect -64 -98 -56 -64
rect -22 -98 -10 -64
rect -64 -124 -10 -98
rect 26 -64 84 -40
rect 26 -98 38 -64
rect 72 -98 84 -64
rect 26 -124 84 -98
rect 120 -64 214 -40
rect 120 -98 132 -64
rect 166 -98 214 -64
rect 120 -124 214 -98
rect 250 -64 352 -40
rect 250 -98 290 -64
rect 324 -98 352 -64
rect 250 -124 352 -98
rect 388 -64 446 -40
rect 388 -98 400 -64
rect 434 -98 446 -64
rect 388 -124 446 -98
rect 482 -64 536 -40
rect 482 -98 494 -64
rect 528 -98 536 -64
rect 482 -124 536 -98
rect 594 -66 648 -40
rect 594 -100 602 -66
rect 636 -100 648 -66
rect 594 -124 648 -100
rect 684 -64 746 -40
rect 684 -98 696 -64
rect 734 -98 746 -64
rect 684 -124 746 -98
rect 782 -64 836 -40
rect 782 -98 794 -64
rect 828 -98 836 -64
rect 782 -124 836 -98
<< pdiff >>
rect -64 286 -10 310
rect -64 252 -56 286
rect -22 252 -10 286
rect -64 226 -10 252
rect 26 226 84 310
rect 120 286 214 310
rect 120 252 132 286
rect 166 252 214 286
rect 120 226 214 252
rect 250 226 352 310
rect 388 286 442 310
rect 388 252 400 286
rect 434 252 442 286
rect 388 226 442 252
rect 604 286 658 310
rect 604 252 612 286
rect 646 252 658 286
rect 604 226 658 252
rect 694 286 752 310
rect 694 252 706 286
rect 740 252 752 286
rect 694 226 752 252
rect 788 286 850 310
rect 788 252 800 286
rect 838 252 850 286
rect 788 226 850 252
<< ndiffc >>
rect -56 -98 -22 -64
rect 38 -98 72 -64
rect 132 -98 166 -64
rect 290 -98 324 -64
rect 400 -98 434 -64
rect 494 -98 528 -64
rect 602 -100 636 -66
rect 696 -98 734 -64
rect 794 -98 828 -64
<< pdiffc >>
rect -56 252 -22 286
rect 132 252 166 286
rect 400 252 434 286
rect 612 252 646 286
rect 706 252 740 286
rect 800 252 838 286
<< psubdiff >>
rect 890 -64 944 -40
rect 890 -98 900 -64
rect 934 -98 944 -64
rect 890 -124 944 -98
<< nsubdiff >>
rect 496 284 550 308
rect 496 250 506 284
rect 540 250 550 284
rect 496 224 550 250
<< psubdiffcont >>
rect 900 -98 934 -64
<< nsubdiffcont >>
rect 506 250 540 284
<< poly >>
rect -10 310 26 336
rect 84 310 120 336
rect 214 310 250 336
rect 352 310 388 336
rect 658 310 694 336
rect 752 310 788 336
rect -10 202 26 226
rect -116 172 26 202
rect 84 202 120 226
rect 84 200 124 202
rect 84 192 136 200
rect 84 174 162 192
rect 84 172 112 174
rect -116 -48 -80 172
rect 94 170 112 172
rect 100 140 112 170
rect 146 140 162 174
rect -10 112 52 130
rect -10 78 2 112
rect 36 78 52 112
rect -10 60 52 78
rect 100 124 162 140
rect -10 -40 26 60
rect 100 58 136 124
rect 214 80 250 226
rect 352 124 388 226
rect 658 210 694 226
rect 752 210 788 226
rect 446 180 788 210
rect 94 18 136 58
rect 84 -16 136 18
rect 196 62 250 80
rect 196 28 206 62
rect 240 28 250 62
rect 350 106 404 124
rect 350 72 360 106
rect 394 72 404 106
rect 350 54 404 72
rect 446 56 482 180
rect 744 102 798 120
rect 744 68 754 102
rect 788 68 798 102
rect 196 12 250 28
rect 84 -40 120 -16
rect 214 -40 250 12
rect 446 46 516 56
rect 446 12 462 46
rect 496 12 516 46
rect 446 2 516 12
rect 648 46 702 64
rect 744 50 798 68
rect 648 12 658 46
rect 692 12 702 46
rect 352 -40 388 -14
rect 446 -40 482 2
rect 648 -6 702 12
rect 648 -40 684 -6
rect 746 -40 782 50
rect -150 -66 -80 -48
rect -150 -100 -140 -66
rect -106 -100 -80 -66
rect -150 -114 -80 -100
rect -150 -116 -98 -114
rect -10 -192 26 -124
rect 84 -150 120 -124
rect 214 -150 250 -124
rect 352 -192 388 -124
rect 446 -150 482 -124
rect 648 -150 684 -124
rect 746 -150 782 -124
rect -10 -222 388 -192
<< polycont >>
rect 112 140 146 174
rect 2 78 36 112
rect 206 28 240 62
rect 360 72 394 106
rect 754 68 788 102
rect 462 12 496 46
rect 658 12 692 46
rect -140 -100 -106 -66
<< locali >>
rect -115 344 -84 378
rect -50 344 36 378
rect 70 344 218 378
rect 252 344 426 378
rect 460 344 602 378
rect 636 344 756 378
rect 790 344 818 378
rect 134 310 168 344
rect -64 286 -10 310
rect -64 260 -56 286
rect -78 252 -56 260
rect -22 252 -10 286
rect -78 226 -10 252
rect 120 286 178 310
rect 120 252 132 286
rect 166 252 178 286
rect 120 226 178 252
rect 388 286 442 310
rect 510 308 544 344
rect 710 310 746 344
rect 388 252 400 286
rect 434 252 442 286
rect 388 226 442 252
rect -78 28 -44 226
rect 408 192 442 226
rect 496 284 550 308
rect 496 250 506 284
rect 540 250 550 284
rect 496 224 550 250
rect 604 286 658 310
rect 604 252 612 286
rect 646 252 658 286
rect 604 226 658 252
rect 694 286 752 310
rect 694 252 706 286
rect 740 252 752 286
rect 694 226 752 252
rect 788 286 850 310
rect 788 252 800 286
rect 838 262 850 286
rect 838 252 870 262
rect 788 226 870 252
rect 604 198 638 226
rect 100 174 442 192
rect 584 190 638 198
rect 100 140 112 174
rect 146 158 442 174
rect 146 140 162 158
rect -10 112 52 130
rect 100 124 162 140
rect -10 78 2 112
rect 36 78 52 112
rect -10 62 52 78
rect 196 62 248 80
rect 196 28 206 62
rect 240 28 248 62
rect -78 -6 248 28
rect 40 -40 74 -6
rect 282 -40 316 158
rect 574 156 638 190
rect 574 124 608 156
rect 350 106 608 124
rect 350 72 360 106
rect 394 90 608 106
rect 394 72 404 90
rect 350 56 404 72
rect 446 46 516 56
rect 446 12 462 46
rect 496 12 516 46
rect 446 2 516 12
rect 574 -40 608 90
rect 744 102 798 120
rect 744 68 754 102
rect 788 68 798 102
rect 648 46 702 64
rect 744 62 798 68
rect 744 50 788 62
rect 648 12 658 46
rect 692 12 702 46
rect 836 28 870 226
rect 824 26 870 28
rect 648 -6 702 12
rect 822 -4 870 26
rect 812 -8 870 -4
rect 812 -40 856 -8
rect -150 -66 -98 -48
rect -150 -100 -140 -66
rect -106 -100 -98 -66
rect -150 -116 -98 -100
rect -132 -226 -98 -116
rect -64 -64 -10 -40
rect -64 -98 -56 -64
rect -22 -98 -10 -64
rect -64 -124 -10 -98
rect 26 -64 84 -40
rect 26 -98 38 -64
rect 72 -98 84 -64
rect 26 -124 84 -98
rect 120 -48 154 -40
rect 120 -64 178 -48
rect 120 -98 132 -64
rect 166 -98 178 -64
rect 120 -124 178 -98
rect 278 -64 336 -40
rect 278 -98 290 -64
rect 324 -98 336 -64
rect 278 -124 336 -98
rect 388 -64 446 -40
rect 388 -98 400 -64
rect 434 -98 446 -64
rect 388 -124 446 -98
rect 482 -64 536 -40
rect 482 -98 494 -64
rect 528 -98 536 -64
rect 574 -66 648 -40
rect 574 -80 602 -66
rect 482 -124 536 -98
rect 594 -100 602 -80
rect 636 -100 648 -66
rect 594 -124 648 -100
rect 684 -64 746 -40
rect 684 -98 696 -64
rect 734 -98 746 -64
rect 684 -124 746 -98
rect 782 -64 856 -40
rect 782 -98 794 -64
rect 828 -74 856 -64
rect 890 -64 944 -48
rect 828 -98 836 -74
rect 782 -124 836 -98
rect -64 -158 -30 -124
rect 134 -158 168 -124
rect 408 -158 442 -124
rect -64 -192 442 -158
rect 502 -158 536 -124
rect 702 -158 736 -124
rect 502 -192 736 -158
rect 802 -226 836 -124
rect -132 -260 836 -226
rect 890 -98 900 -64
rect 934 -98 944 -64
rect 890 -114 944 -98
rect 890 -238 924 -114
<< viali >>
rect -84 344 -50 378
rect 36 344 70 378
rect 218 344 252 378
rect 426 344 460 378
rect 602 344 636 378
rect 756 344 790 378
rect 400 -98 434 -64
rect 890 -272 924 -238
<< metal1 >>
rect -186 378 976 388
rect -186 344 -84 378
rect -50 344 36 378
rect 70 344 218 378
rect 252 344 426 378
rect 460 344 602 378
rect 636 344 756 378
rect 790 344 976 378
rect -186 338 976 344
rect 388 -64 446 -52
rect 388 -98 400 -64
rect 434 -98 446 -64
rect 388 -232 446 -98
rect -186 -238 976 -232
rect -186 -272 890 -238
rect 924 -272 976 -238
rect -186 -282 976 -272
<< labels >>
rlabel metal1 -186 362 -186 362 7 VDD
rlabel metal1 -186 -260 -186 -260 7 GND
rlabel locali 516 28 516 28 3 clk
rlabel locali 196 32 196 32 7 out
rlabel locali 20 130 20 130 1 clkbar
rlabel locali 772 120 772 120 1 vinp
rlabel locali 674 64 674 64 1 vinm
<< end >>
