magic
tech minimum
timestamp 0
<< end >>
