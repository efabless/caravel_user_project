magic
tech sky130A
timestamp 1641072977
<< nwell >>
rect -88 552 1192 644
rect -88 248 4 552
rect 261 438 345 552
rect 685 437 769 552
rect 1107 438 1191 552
rect -88 214 1 248
rect -86 109 1 214
rect -86 -78 259 109
rect 1260 103 1404 109
rect 1260 89 1443 103
rect 1253 5 1443 89
rect 1272 2 1443 5
rect 1271 -1 1443 2
rect 1271 -78 1412 -1
rect -86 -3816 1 -78
rect 1358 -291 1442 -288
rect 1272 -478 1442 -291
rect 1358 -493 1442 -478
rect 1358 -691 1442 -688
rect 1272 -878 1442 -691
rect 1358 -893 1442 -878
rect 1357 -1091 1441 -1088
rect 1271 -1278 1441 -1091
rect 1357 -1293 1441 -1278
rect 1358 -1491 1442 -1488
rect 1272 -1678 1442 -1491
rect 1358 -1693 1442 -1678
rect 1356 -1891 1440 -1888
rect 1270 -2078 1440 -1891
rect 1356 -2093 1440 -2078
rect 1358 -2291 1442 -2288
rect 1272 -2478 1442 -2291
rect 1358 -2493 1442 -2478
rect 1358 -2691 1442 -2688
rect 1272 -2878 1442 -2691
rect 1358 -2893 1442 -2878
rect 1358 -3091 1442 -3088
rect 1272 -3278 1442 -3091
rect 1358 -3293 1442 -3278
rect 1358 -3491 1442 -3488
rect 1272 -3678 1442 -3491
rect 1358 -3693 1442 -3678
rect -86 -4000 68 -3816
rect -86 -4050 134 -4000
rect -86 -4100 135 -4050
rect 474 -4100 558 -4000
rect 896 -4100 980 -3998
rect -86 -4187 981 -4100
<< nmos >>
rect 1477 -349 1519 -334
rect 1477 -447 1519 -432
rect 1477 -749 1519 -734
rect 1477 -847 1519 -832
rect 1476 -1149 1518 -1134
rect 1476 -1247 1518 -1232
rect 1477 -1549 1519 -1534
rect 1477 -1647 1519 -1632
rect 1475 -1949 1517 -1934
rect 1475 -2047 1517 -2032
rect 1477 -2349 1519 -2334
rect 1477 -2447 1519 -2432
rect 1477 -2749 1519 -2734
rect 1477 -2847 1519 -2832
rect 1477 -3149 1519 -3134
rect 1477 -3247 1519 -3232
rect 1477 -3549 1519 -3534
rect 1477 -3647 1519 -3632
<< pmos >>
rect 1382 -349 1424 -334
rect 1382 -447 1424 -432
rect 1382 -749 1424 -734
rect 1382 -847 1424 -832
rect 1381 -1149 1423 -1134
rect 1381 -1247 1423 -1232
rect 1382 -1549 1424 -1534
rect 1382 -1647 1424 -1632
rect 1380 -1949 1422 -1934
rect 1380 -2047 1422 -2032
rect 1382 -2349 1424 -2334
rect 1382 -2447 1424 -2432
rect 1382 -2749 1424 -2734
rect 1382 -2847 1424 -2832
rect 1382 -3149 1424 -3134
rect 1382 -3247 1424 -3232
rect 1382 -3549 1424 -3534
rect 1382 -3647 1424 -3632
<< ndiff >>
rect 1477 -311 1519 -306
rect 1477 -328 1490 -311
rect 1507 -328 1519 -311
rect 1477 -334 1519 -328
rect 1477 -355 1519 -349
rect 1477 -372 1490 -355
rect 1507 -372 1519 -355
rect 1477 -377 1519 -372
rect 1477 -409 1519 -404
rect 1477 -426 1490 -409
rect 1507 -426 1519 -409
rect 1477 -432 1519 -426
rect 1477 -453 1519 -447
rect 1477 -470 1490 -453
rect 1507 -470 1519 -453
rect 1477 -475 1519 -470
rect 1477 -711 1519 -706
rect 1477 -728 1490 -711
rect 1507 -728 1519 -711
rect 1477 -734 1519 -728
rect 1477 -755 1519 -749
rect 1477 -772 1490 -755
rect 1507 -772 1519 -755
rect 1477 -777 1519 -772
rect 1477 -809 1519 -804
rect 1477 -826 1490 -809
rect 1507 -826 1519 -809
rect 1477 -832 1519 -826
rect 1477 -853 1519 -847
rect 1477 -870 1490 -853
rect 1507 -870 1519 -853
rect 1477 -875 1519 -870
rect 1476 -1111 1518 -1106
rect 1476 -1128 1489 -1111
rect 1506 -1128 1518 -1111
rect 1476 -1134 1518 -1128
rect 1476 -1155 1518 -1149
rect 1476 -1172 1489 -1155
rect 1506 -1172 1518 -1155
rect 1476 -1177 1518 -1172
rect 1476 -1209 1518 -1204
rect 1476 -1226 1489 -1209
rect 1506 -1226 1518 -1209
rect 1476 -1232 1518 -1226
rect 1476 -1253 1518 -1247
rect 1476 -1270 1489 -1253
rect 1506 -1270 1518 -1253
rect 1476 -1275 1518 -1270
rect 1477 -1511 1519 -1506
rect 1477 -1528 1490 -1511
rect 1507 -1528 1519 -1511
rect 1477 -1534 1519 -1528
rect 1477 -1555 1519 -1549
rect 1477 -1572 1490 -1555
rect 1507 -1572 1519 -1555
rect 1477 -1577 1519 -1572
rect 1477 -1609 1519 -1604
rect 1477 -1626 1490 -1609
rect 1507 -1626 1519 -1609
rect 1477 -1632 1519 -1626
rect 1477 -1653 1519 -1647
rect 1477 -1670 1490 -1653
rect 1507 -1670 1519 -1653
rect 1477 -1675 1519 -1670
rect 1475 -1911 1517 -1906
rect 1475 -1928 1488 -1911
rect 1505 -1928 1517 -1911
rect 1475 -1934 1517 -1928
rect 1475 -1955 1517 -1949
rect 1475 -1972 1488 -1955
rect 1505 -1972 1517 -1955
rect 1475 -1977 1517 -1972
rect 1475 -2009 1517 -2004
rect 1475 -2026 1488 -2009
rect 1505 -2026 1517 -2009
rect 1475 -2032 1517 -2026
rect 1475 -2053 1517 -2047
rect 1475 -2070 1488 -2053
rect 1505 -2070 1517 -2053
rect 1475 -2075 1517 -2070
rect 1477 -2311 1519 -2306
rect 1477 -2328 1490 -2311
rect 1507 -2328 1519 -2311
rect 1477 -2334 1519 -2328
rect 1477 -2355 1519 -2349
rect 1477 -2372 1490 -2355
rect 1507 -2372 1519 -2355
rect 1477 -2377 1519 -2372
rect 1477 -2409 1519 -2404
rect 1477 -2426 1490 -2409
rect 1507 -2426 1519 -2409
rect 1477 -2432 1519 -2426
rect 1477 -2453 1519 -2447
rect 1477 -2470 1490 -2453
rect 1507 -2470 1519 -2453
rect 1477 -2475 1519 -2470
rect 1477 -2711 1519 -2706
rect 1477 -2728 1490 -2711
rect 1507 -2728 1519 -2711
rect 1477 -2734 1519 -2728
rect 1477 -2755 1519 -2749
rect 1477 -2772 1490 -2755
rect 1507 -2772 1519 -2755
rect 1477 -2777 1519 -2772
rect 1477 -2809 1519 -2804
rect 1477 -2826 1490 -2809
rect 1507 -2826 1519 -2809
rect 1477 -2832 1519 -2826
rect 1477 -2853 1519 -2847
rect 1477 -2870 1490 -2853
rect 1507 -2870 1519 -2853
rect 1477 -2875 1519 -2870
rect 1477 -3111 1519 -3106
rect 1477 -3128 1490 -3111
rect 1507 -3128 1519 -3111
rect 1477 -3134 1519 -3128
rect 1477 -3155 1519 -3149
rect 1477 -3172 1490 -3155
rect 1507 -3172 1519 -3155
rect 1477 -3177 1519 -3172
rect 1477 -3209 1519 -3204
rect 1477 -3226 1490 -3209
rect 1507 -3226 1519 -3209
rect 1477 -3232 1519 -3226
rect 1477 -3253 1519 -3247
rect 1477 -3270 1490 -3253
rect 1507 -3270 1519 -3253
rect 1477 -3275 1519 -3270
rect 1477 -3511 1519 -3506
rect 1477 -3528 1490 -3511
rect 1507 -3528 1519 -3511
rect 1477 -3534 1519 -3528
rect 1477 -3555 1519 -3549
rect 1477 -3572 1490 -3555
rect 1507 -3572 1519 -3555
rect 1477 -3577 1519 -3572
rect 1477 -3609 1519 -3604
rect 1477 -3626 1490 -3609
rect 1507 -3626 1519 -3609
rect 1477 -3632 1519 -3626
rect 1477 -3653 1519 -3647
rect 1477 -3670 1490 -3653
rect 1507 -3670 1519 -3653
rect 1477 -3675 1519 -3670
<< pdiff >>
rect 1382 -311 1424 -306
rect 1382 -328 1394 -311
rect 1411 -328 1424 -311
rect 1382 -334 1424 -328
rect 1382 -355 1424 -349
rect 1382 -372 1394 -355
rect 1411 -372 1424 -355
rect 1382 -377 1424 -372
rect 1382 -409 1424 -404
rect 1382 -426 1394 -409
rect 1411 -426 1424 -409
rect 1382 -432 1424 -426
rect 1382 -453 1424 -447
rect 1382 -470 1394 -453
rect 1411 -470 1424 -453
rect 1382 -475 1424 -470
rect 1382 -711 1424 -706
rect 1382 -728 1394 -711
rect 1411 -728 1424 -711
rect 1382 -734 1424 -728
rect 1382 -755 1424 -749
rect 1382 -772 1394 -755
rect 1411 -772 1424 -755
rect 1382 -777 1424 -772
rect 1382 -809 1424 -804
rect 1382 -826 1394 -809
rect 1411 -826 1424 -809
rect 1382 -832 1424 -826
rect 1382 -853 1424 -847
rect 1382 -870 1394 -853
rect 1411 -870 1424 -853
rect 1382 -875 1424 -870
rect 1381 -1111 1423 -1106
rect 1381 -1128 1393 -1111
rect 1410 -1128 1423 -1111
rect 1381 -1134 1423 -1128
rect 1381 -1155 1423 -1149
rect 1381 -1172 1393 -1155
rect 1410 -1172 1423 -1155
rect 1381 -1177 1423 -1172
rect 1381 -1209 1423 -1204
rect 1381 -1226 1393 -1209
rect 1410 -1226 1423 -1209
rect 1381 -1232 1423 -1226
rect 1381 -1253 1423 -1247
rect 1381 -1270 1393 -1253
rect 1410 -1270 1423 -1253
rect 1381 -1275 1423 -1270
rect 1382 -1511 1424 -1506
rect 1382 -1528 1394 -1511
rect 1411 -1528 1424 -1511
rect 1382 -1534 1424 -1528
rect 1382 -1555 1424 -1549
rect 1382 -1572 1394 -1555
rect 1411 -1572 1424 -1555
rect 1382 -1577 1424 -1572
rect 1382 -1609 1424 -1604
rect 1382 -1626 1394 -1609
rect 1411 -1626 1424 -1609
rect 1382 -1632 1424 -1626
rect 1382 -1653 1424 -1647
rect 1382 -1670 1394 -1653
rect 1411 -1670 1424 -1653
rect 1382 -1675 1424 -1670
rect 1380 -1911 1422 -1906
rect 1380 -1928 1392 -1911
rect 1409 -1928 1422 -1911
rect 1380 -1934 1422 -1928
rect 1380 -1955 1422 -1949
rect 1380 -1972 1392 -1955
rect 1409 -1972 1422 -1955
rect 1380 -1977 1422 -1972
rect 1380 -2009 1422 -2004
rect 1380 -2026 1392 -2009
rect 1409 -2026 1422 -2009
rect 1380 -2032 1422 -2026
rect 1380 -2053 1422 -2047
rect 1380 -2070 1392 -2053
rect 1409 -2070 1422 -2053
rect 1380 -2075 1422 -2070
rect 1382 -2311 1424 -2306
rect 1382 -2328 1394 -2311
rect 1411 -2328 1424 -2311
rect 1382 -2334 1424 -2328
rect 1382 -2355 1424 -2349
rect 1382 -2372 1394 -2355
rect 1411 -2372 1424 -2355
rect 1382 -2377 1424 -2372
rect 1382 -2409 1424 -2404
rect 1382 -2426 1394 -2409
rect 1411 -2426 1424 -2409
rect 1382 -2432 1424 -2426
rect 1382 -2453 1424 -2447
rect 1382 -2470 1394 -2453
rect 1411 -2470 1424 -2453
rect 1382 -2475 1424 -2470
rect 1382 -2711 1424 -2706
rect 1382 -2728 1394 -2711
rect 1411 -2728 1424 -2711
rect 1382 -2734 1424 -2728
rect 1382 -2755 1424 -2749
rect 1382 -2772 1394 -2755
rect 1411 -2772 1424 -2755
rect 1382 -2777 1424 -2772
rect 1382 -2809 1424 -2804
rect 1382 -2826 1394 -2809
rect 1411 -2826 1424 -2809
rect 1382 -2832 1424 -2826
rect 1382 -2853 1424 -2847
rect 1382 -2870 1394 -2853
rect 1411 -2870 1424 -2853
rect 1382 -2875 1424 -2870
rect 1382 -3111 1424 -3106
rect 1382 -3128 1394 -3111
rect 1411 -3128 1424 -3111
rect 1382 -3134 1424 -3128
rect 1382 -3155 1424 -3149
rect 1382 -3172 1394 -3155
rect 1411 -3172 1424 -3155
rect 1382 -3177 1424 -3172
rect 1382 -3209 1424 -3204
rect 1382 -3226 1394 -3209
rect 1411 -3226 1424 -3209
rect 1382 -3232 1424 -3226
rect 1382 -3253 1424 -3247
rect 1382 -3270 1394 -3253
rect 1411 -3270 1424 -3253
rect 1382 -3275 1424 -3270
rect 1382 -3511 1424 -3506
rect 1382 -3528 1394 -3511
rect 1411 -3528 1424 -3511
rect 1382 -3534 1424 -3528
rect 1382 -3555 1424 -3549
rect 1382 -3572 1394 -3555
rect 1411 -3572 1424 -3555
rect 1382 -3577 1424 -3572
rect 1382 -3609 1424 -3604
rect 1382 -3626 1394 -3609
rect 1411 -3626 1424 -3609
rect 1382 -3632 1424 -3626
rect 1382 -3653 1424 -3647
rect 1382 -3670 1394 -3653
rect 1411 -3670 1424 -3653
rect 1382 -3675 1424 -3670
<< ndiffc >>
rect 1490 -328 1507 -311
rect 1490 -372 1507 -355
rect 1490 -426 1507 -409
rect 1490 -470 1507 -453
rect 1490 -728 1507 -711
rect 1490 -772 1507 -755
rect 1490 -826 1507 -809
rect 1490 -870 1507 -853
rect 1489 -1128 1506 -1111
rect 1489 -1172 1506 -1155
rect 1489 -1226 1506 -1209
rect 1489 -1270 1506 -1253
rect 1490 -1528 1507 -1511
rect 1490 -1572 1507 -1555
rect 1490 -1626 1507 -1609
rect 1490 -1670 1507 -1653
rect 1488 -1928 1505 -1911
rect 1488 -1972 1505 -1955
rect 1488 -2026 1505 -2009
rect 1488 -2070 1505 -2053
rect 1490 -2328 1507 -2311
rect 1490 -2372 1507 -2355
rect 1490 -2426 1507 -2409
rect 1490 -2470 1507 -2453
rect 1490 -2728 1507 -2711
rect 1490 -2772 1507 -2755
rect 1490 -2826 1507 -2809
rect 1490 -2870 1507 -2853
rect 1490 -3128 1507 -3111
rect 1490 -3172 1507 -3155
rect 1490 -3226 1507 -3209
rect 1490 -3270 1507 -3253
rect 1490 -3528 1507 -3511
rect 1490 -3572 1507 -3555
rect 1490 -3626 1507 -3609
rect 1490 -3670 1507 -3653
<< pdiffc >>
rect 1394 -328 1411 -311
rect 1394 -372 1411 -355
rect 1394 -426 1411 -409
rect 1394 -470 1411 -453
rect 1394 -728 1411 -711
rect 1394 -772 1411 -755
rect 1394 -826 1411 -809
rect 1394 -870 1411 -853
rect 1393 -1128 1410 -1111
rect 1393 -1172 1410 -1155
rect 1393 -1226 1410 -1209
rect 1393 -1270 1410 -1253
rect 1394 -1528 1411 -1511
rect 1394 -1572 1411 -1555
rect 1394 -1626 1411 -1609
rect 1394 -1670 1411 -1653
rect 1392 -1928 1409 -1911
rect 1392 -1972 1409 -1955
rect 1392 -2026 1409 -2009
rect 1392 -2070 1409 -2053
rect 1394 -2328 1411 -2311
rect 1394 -2372 1411 -2355
rect 1394 -2426 1411 -2409
rect 1394 -2470 1411 -2453
rect 1394 -2728 1411 -2711
rect 1394 -2772 1411 -2755
rect 1394 -2826 1411 -2809
rect 1394 -2870 1411 -2853
rect 1394 -3128 1411 -3111
rect 1394 -3172 1411 -3155
rect 1394 -3226 1411 -3209
rect 1394 -3270 1411 -3253
rect 1394 -3528 1411 -3511
rect 1394 -3572 1411 -3555
rect 1394 -3626 1411 -3609
rect 1394 -3670 1411 -3653
<< poly >>
rect 1331 -332 1374 -322
rect 1331 -351 1336 -332
rect 1353 -334 1374 -332
rect 1527 -332 1563 -322
rect 1527 -334 1541 -332
rect 1353 -349 1382 -334
rect 1424 -349 1477 -334
rect 1519 -349 1541 -334
rect 1353 -351 1374 -349
rect 1331 -361 1374 -351
rect 1527 -351 1541 -349
rect 1558 -351 1563 -332
rect 1527 -361 1563 -351
rect 1331 -430 1374 -420
rect 1331 -449 1336 -430
rect 1353 -432 1374 -430
rect 1527 -430 1563 -420
rect 1527 -432 1541 -430
rect 1353 -447 1382 -432
rect 1424 -447 1477 -432
rect 1519 -447 1541 -432
rect 1353 -449 1374 -447
rect 1331 -459 1374 -449
rect 1527 -449 1541 -447
rect 1558 -449 1563 -430
rect 1527 -459 1563 -449
rect 1331 -732 1374 -722
rect 1331 -751 1336 -732
rect 1353 -734 1374 -732
rect 1527 -732 1563 -722
rect 1527 -734 1541 -732
rect 1353 -749 1382 -734
rect 1424 -749 1477 -734
rect 1519 -749 1541 -734
rect 1353 -751 1374 -749
rect 1331 -761 1374 -751
rect 1527 -751 1541 -749
rect 1558 -751 1563 -732
rect 1527 -761 1563 -751
rect 1331 -830 1374 -820
rect 1331 -849 1336 -830
rect 1353 -832 1374 -830
rect 1527 -830 1563 -820
rect 1527 -832 1541 -830
rect 1353 -847 1382 -832
rect 1424 -847 1477 -832
rect 1519 -847 1541 -832
rect 1353 -849 1374 -847
rect 1331 -859 1374 -849
rect 1527 -849 1541 -847
rect 1558 -849 1563 -830
rect 1527 -859 1563 -849
rect 1330 -1132 1373 -1122
rect 1330 -1151 1335 -1132
rect 1352 -1134 1373 -1132
rect 1526 -1132 1562 -1122
rect 1526 -1134 1540 -1132
rect 1352 -1149 1381 -1134
rect 1423 -1149 1476 -1134
rect 1518 -1149 1540 -1134
rect 1352 -1151 1373 -1149
rect 1330 -1161 1373 -1151
rect 1526 -1151 1540 -1149
rect 1557 -1151 1562 -1132
rect 1526 -1161 1562 -1151
rect 1330 -1230 1373 -1220
rect 1330 -1249 1335 -1230
rect 1352 -1232 1373 -1230
rect 1526 -1230 1562 -1220
rect 1526 -1232 1540 -1230
rect 1352 -1247 1381 -1232
rect 1423 -1247 1476 -1232
rect 1518 -1247 1540 -1232
rect 1352 -1249 1373 -1247
rect 1330 -1259 1373 -1249
rect 1526 -1249 1540 -1247
rect 1557 -1249 1562 -1230
rect 1526 -1259 1562 -1249
rect 1331 -1532 1374 -1522
rect 1331 -1551 1336 -1532
rect 1353 -1534 1374 -1532
rect 1527 -1532 1563 -1522
rect 1527 -1534 1541 -1532
rect 1353 -1549 1382 -1534
rect 1424 -1549 1477 -1534
rect 1519 -1549 1541 -1534
rect 1353 -1551 1374 -1549
rect 1331 -1561 1374 -1551
rect 1527 -1551 1541 -1549
rect 1558 -1551 1563 -1532
rect 1527 -1561 1563 -1551
rect 1331 -1630 1374 -1620
rect 1331 -1649 1336 -1630
rect 1353 -1632 1374 -1630
rect 1527 -1630 1563 -1620
rect 1527 -1632 1541 -1630
rect 1353 -1647 1382 -1632
rect 1424 -1647 1477 -1632
rect 1519 -1647 1541 -1632
rect 1353 -1649 1374 -1647
rect 1331 -1659 1374 -1649
rect 1527 -1649 1541 -1647
rect 1558 -1649 1563 -1630
rect 1527 -1659 1563 -1649
rect 1329 -1932 1372 -1922
rect 1329 -1951 1334 -1932
rect 1351 -1934 1372 -1932
rect 1525 -1932 1561 -1922
rect 1525 -1934 1539 -1932
rect 1351 -1949 1380 -1934
rect 1422 -1949 1475 -1934
rect 1517 -1949 1539 -1934
rect 1351 -1951 1372 -1949
rect 1329 -1961 1372 -1951
rect 1525 -1951 1539 -1949
rect 1556 -1951 1561 -1932
rect 1525 -1961 1561 -1951
rect 1329 -2030 1372 -2020
rect 1329 -2049 1334 -2030
rect 1351 -2032 1372 -2030
rect 1525 -2030 1561 -2020
rect 1525 -2032 1539 -2030
rect 1351 -2047 1380 -2032
rect 1422 -2047 1475 -2032
rect 1517 -2047 1539 -2032
rect 1351 -2049 1372 -2047
rect 1329 -2059 1372 -2049
rect 1525 -2049 1539 -2047
rect 1556 -2049 1561 -2030
rect 1525 -2059 1561 -2049
rect 1331 -2332 1374 -2322
rect 1331 -2351 1336 -2332
rect 1353 -2334 1374 -2332
rect 1527 -2332 1563 -2322
rect 1527 -2334 1541 -2332
rect 1353 -2349 1382 -2334
rect 1424 -2349 1477 -2334
rect 1519 -2349 1541 -2334
rect 1353 -2351 1374 -2349
rect 1331 -2361 1374 -2351
rect 1527 -2351 1541 -2349
rect 1558 -2351 1563 -2332
rect 1527 -2361 1563 -2351
rect 1331 -2430 1374 -2420
rect 1331 -2449 1336 -2430
rect 1353 -2432 1374 -2430
rect 1527 -2430 1563 -2420
rect 1527 -2432 1541 -2430
rect 1353 -2447 1382 -2432
rect 1424 -2447 1477 -2432
rect 1519 -2447 1541 -2432
rect 1353 -2449 1374 -2447
rect 1331 -2459 1374 -2449
rect 1527 -2449 1541 -2447
rect 1558 -2449 1563 -2430
rect 1527 -2459 1563 -2449
rect 1331 -2732 1374 -2722
rect 1331 -2751 1336 -2732
rect 1353 -2734 1374 -2732
rect 1527 -2732 1563 -2722
rect 1527 -2734 1541 -2732
rect 1353 -2749 1382 -2734
rect 1424 -2749 1477 -2734
rect 1519 -2749 1541 -2734
rect 1353 -2751 1374 -2749
rect 1331 -2761 1374 -2751
rect 1527 -2751 1541 -2749
rect 1558 -2751 1563 -2732
rect 1527 -2761 1563 -2751
rect 1331 -2830 1374 -2820
rect 1331 -2849 1336 -2830
rect 1353 -2832 1374 -2830
rect 1527 -2830 1563 -2820
rect 1527 -2832 1541 -2830
rect 1353 -2847 1382 -2832
rect 1424 -2847 1477 -2832
rect 1519 -2847 1541 -2832
rect 1353 -2849 1374 -2847
rect 1331 -2859 1374 -2849
rect 1527 -2849 1541 -2847
rect 1558 -2849 1563 -2830
rect 1527 -2859 1563 -2849
rect 1331 -3132 1374 -3122
rect 1331 -3151 1336 -3132
rect 1353 -3134 1374 -3132
rect 1527 -3132 1563 -3122
rect 1527 -3134 1541 -3132
rect 1353 -3149 1382 -3134
rect 1424 -3149 1477 -3134
rect 1519 -3149 1541 -3134
rect 1353 -3151 1374 -3149
rect 1331 -3161 1374 -3151
rect 1527 -3151 1541 -3149
rect 1558 -3151 1563 -3132
rect 1527 -3161 1563 -3151
rect 1331 -3230 1374 -3220
rect 1331 -3249 1336 -3230
rect 1353 -3232 1374 -3230
rect 1527 -3230 1563 -3220
rect 1527 -3232 1541 -3230
rect 1353 -3247 1382 -3232
rect 1424 -3247 1477 -3232
rect 1519 -3247 1541 -3232
rect 1353 -3249 1374 -3247
rect 1331 -3259 1374 -3249
rect 1527 -3249 1541 -3247
rect 1558 -3249 1563 -3230
rect 1527 -3259 1563 -3249
rect 1331 -3532 1374 -3522
rect 1331 -3551 1336 -3532
rect 1353 -3534 1374 -3532
rect 1527 -3532 1563 -3522
rect 1527 -3534 1541 -3532
rect 1353 -3549 1382 -3534
rect 1424 -3549 1477 -3534
rect 1519 -3549 1541 -3534
rect 1353 -3551 1374 -3549
rect 1331 -3561 1374 -3551
rect 1527 -3551 1541 -3549
rect 1558 -3551 1563 -3532
rect 1527 -3561 1563 -3551
rect 1331 -3630 1374 -3620
rect 1331 -3649 1336 -3630
rect 1353 -3632 1374 -3630
rect 1527 -3630 1563 -3620
rect 1527 -3632 1541 -3630
rect 1353 -3647 1382 -3632
rect 1424 -3647 1477 -3632
rect 1519 -3647 1541 -3632
rect 1353 -3649 1374 -3647
rect 1331 -3659 1374 -3649
rect 1527 -3649 1541 -3647
rect 1558 -3649 1563 -3630
rect 1527 -3659 1563 -3649
<< polycont >>
rect 1336 -351 1353 -332
rect 1541 -351 1558 -332
rect 1336 -449 1353 -430
rect 1541 -449 1558 -430
rect 1336 -751 1353 -732
rect 1541 -751 1558 -732
rect 1336 -849 1353 -830
rect 1541 -849 1558 -830
rect 1335 -1151 1352 -1132
rect 1540 -1151 1557 -1132
rect 1335 -1249 1352 -1230
rect 1540 -1249 1557 -1230
rect 1336 -1551 1353 -1532
rect 1541 -1551 1558 -1532
rect 1336 -1649 1353 -1630
rect 1541 -1649 1558 -1630
rect 1334 -1951 1351 -1932
rect 1539 -1951 1556 -1932
rect 1334 -2049 1351 -2030
rect 1539 -2049 1556 -2030
rect 1336 -2351 1353 -2332
rect 1541 -2351 1558 -2332
rect 1336 -2449 1353 -2430
rect 1541 -2449 1558 -2430
rect 1336 -2751 1353 -2732
rect 1541 -2751 1558 -2732
rect 1336 -2849 1353 -2830
rect 1541 -2849 1558 -2830
rect 1336 -3151 1353 -3132
rect 1541 -3151 1558 -3132
rect 1336 -3249 1353 -3230
rect 1541 -3249 1558 -3230
rect 1336 -3551 1353 -3532
rect 1541 -3551 1558 -3532
rect 1336 -3649 1353 -3630
rect 1541 -3649 1558 -3630
<< locali >>
rect 235 289 255 360
rect 659 293 679 357
rect 235 224 264 289
rect 235 204 291 224
rect 337 196 364 277
rect 659 202 690 293
rect 761 202 788 274
rect 1081 229 1108 304
rect 1192 280 1212 281
rect 1081 202 1147 229
rect 1189 223 1212 280
rect 1192 216 1212 223
rect 1443 -306 1463 -295
rect 1382 -311 1519 -306
rect 1331 -332 1365 -322
rect 1382 -328 1394 -311
rect 1411 -326 1490 -311
rect 1411 -328 1424 -326
rect 1382 -332 1424 -328
rect 1477 -328 1490 -326
rect 1507 -328 1519 -311
rect 1477 -332 1519 -328
rect 1536 -332 1563 -322
rect 1331 -351 1336 -332
rect 1353 -351 1365 -332
rect 1536 -351 1541 -332
rect 1558 -351 1563 -332
rect 1331 -361 1365 -351
rect 1382 -355 1424 -351
rect 1382 -372 1394 -355
rect 1411 -372 1424 -355
rect 1382 -377 1424 -372
rect 1477 -355 1519 -351
rect 1477 -372 1490 -355
rect 1507 -372 1519 -355
rect 1536 -361 1563 -351
rect 1477 -377 1519 -372
rect 1392 -404 1411 -377
rect 1490 -404 1509 -377
rect 1382 -409 1424 -404
rect 1331 -430 1365 -420
rect 1382 -426 1394 -409
rect 1411 -426 1424 -409
rect 1382 -430 1424 -426
rect 1477 -409 1519 -404
rect 1477 -426 1490 -409
rect 1507 -426 1519 -409
rect 1477 -430 1519 -426
rect 1536 -430 1563 -420
rect 1331 -449 1336 -430
rect 1353 -449 1365 -430
rect 1536 -449 1541 -430
rect 1558 -449 1563 -430
rect 1331 -459 1365 -449
rect 1382 -453 1424 -449
rect 1382 -470 1394 -453
rect 1411 -455 1424 -453
rect 1477 -453 1519 -449
rect 1477 -455 1490 -453
rect 1411 -470 1490 -455
rect 1507 -470 1519 -453
rect 1536 -459 1563 -449
rect 1382 -475 1519 -470
rect 1443 -486 1463 -475
rect 1443 -706 1463 -695
rect 1382 -711 1519 -706
rect 1331 -732 1365 -722
rect 1382 -728 1394 -711
rect 1411 -726 1490 -711
rect 1411 -728 1424 -726
rect 1382 -732 1424 -728
rect 1477 -728 1490 -726
rect 1507 -728 1519 -711
rect 1477 -732 1519 -728
rect 1536 -732 1563 -722
rect 1331 -751 1336 -732
rect 1353 -751 1365 -732
rect 1536 -751 1541 -732
rect 1558 -751 1563 -732
rect 1331 -761 1365 -751
rect 1382 -755 1424 -751
rect 1382 -772 1394 -755
rect 1411 -772 1424 -755
rect 1382 -777 1424 -772
rect 1477 -755 1519 -751
rect 1477 -772 1490 -755
rect 1507 -772 1519 -755
rect 1536 -761 1563 -751
rect 1477 -777 1519 -772
rect 1392 -804 1411 -777
rect 1490 -804 1509 -777
rect 1382 -809 1424 -804
rect 1331 -830 1365 -820
rect 1382 -826 1394 -809
rect 1411 -826 1424 -809
rect 1382 -830 1424 -826
rect 1477 -809 1519 -804
rect 1477 -826 1490 -809
rect 1507 -826 1519 -809
rect 1477 -830 1519 -826
rect 1536 -830 1563 -820
rect 1331 -849 1336 -830
rect 1353 -849 1365 -830
rect 1536 -849 1541 -830
rect 1558 -849 1563 -830
rect 1331 -859 1365 -849
rect 1382 -853 1424 -849
rect 1382 -870 1394 -853
rect 1411 -855 1424 -853
rect 1477 -853 1519 -849
rect 1477 -855 1490 -853
rect 1411 -870 1490 -855
rect 1507 -870 1519 -853
rect 1536 -859 1563 -849
rect 1382 -875 1519 -870
rect 1443 -886 1463 -875
rect 1442 -1106 1462 -1095
rect 1381 -1111 1518 -1106
rect 1330 -1132 1364 -1122
rect 1381 -1128 1393 -1111
rect 1410 -1126 1489 -1111
rect 1410 -1128 1423 -1126
rect 1381 -1132 1423 -1128
rect 1476 -1128 1489 -1126
rect 1506 -1128 1518 -1111
rect 1476 -1132 1518 -1128
rect 1535 -1132 1562 -1122
rect 1330 -1151 1335 -1132
rect 1352 -1151 1364 -1132
rect 1535 -1151 1540 -1132
rect 1557 -1151 1562 -1132
rect 1330 -1161 1364 -1151
rect 1381 -1155 1423 -1151
rect 1381 -1172 1393 -1155
rect 1410 -1172 1423 -1155
rect 1381 -1177 1423 -1172
rect 1476 -1155 1518 -1151
rect 1476 -1172 1489 -1155
rect 1506 -1172 1518 -1155
rect 1535 -1161 1562 -1151
rect 1476 -1177 1518 -1172
rect 1391 -1204 1410 -1177
rect 1489 -1204 1508 -1177
rect 1381 -1209 1423 -1204
rect 1330 -1230 1364 -1220
rect 1381 -1226 1393 -1209
rect 1410 -1226 1423 -1209
rect 1381 -1230 1423 -1226
rect 1476 -1209 1518 -1204
rect 1476 -1226 1489 -1209
rect 1506 -1226 1518 -1209
rect 1476 -1230 1518 -1226
rect 1535 -1230 1562 -1220
rect 1330 -1249 1335 -1230
rect 1352 -1249 1364 -1230
rect 1535 -1249 1540 -1230
rect 1557 -1249 1562 -1230
rect 1330 -1259 1364 -1249
rect 1381 -1253 1423 -1249
rect 1381 -1270 1393 -1253
rect 1410 -1255 1423 -1253
rect 1476 -1253 1518 -1249
rect 1476 -1255 1489 -1253
rect 1410 -1270 1489 -1255
rect 1506 -1270 1518 -1253
rect 1535 -1259 1562 -1249
rect 1381 -1275 1518 -1270
rect 1442 -1286 1462 -1275
rect 1443 -1506 1463 -1495
rect 1382 -1511 1519 -1506
rect 1331 -1532 1365 -1522
rect 1382 -1528 1394 -1511
rect 1411 -1526 1490 -1511
rect 1411 -1528 1424 -1526
rect 1382 -1532 1424 -1528
rect 1477 -1528 1490 -1526
rect 1507 -1528 1519 -1511
rect 1477 -1532 1519 -1528
rect 1536 -1532 1563 -1522
rect 1331 -1551 1336 -1532
rect 1353 -1551 1365 -1532
rect 1536 -1551 1541 -1532
rect 1558 -1551 1563 -1532
rect 1331 -1561 1365 -1551
rect 1382 -1555 1424 -1551
rect 1382 -1572 1394 -1555
rect 1411 -1572 1424 -1555
rect 1382 -1577 1424 -1572
rect 1477 -1555 1519 -1551
rect 1477 -1572 1490 -1555
rect 1507 -1572 1519 -1555
rect 1536 -1561 1563 -1551
rect 1477 -1577 1519 -1572
rect 1392 -1604 1411 -1577
rect 1490 -1604 1509 -1577
rect 1382 -1609 1424 -1604
rect 1331 -1630 1365 -1620
rect 1382 -1626 1394 -1609
rect 1411 -1626 1424 -1609
rect 1382 -1630 1424 -1626
rect 1477 -1609 1519 -1604
rect 1477 -1626 1490 -1609
rect 1507 -1626 1519 -1609
rect 1477 -1630 1519 -1626
rect 1536 -1630 1563 -1620
rect 1331 -1649 1336 -1630
rect 1353 -1649 1365 -1630
rect 1536 -1649 1541 -1630
rect 1558 -1649 1563 -1630
rect 1331 -1659 1365 -1649
rect 1382 -1653 1424 -1649
rect 1382 -1670 1394 -1653
rect 1411 -1655 1424 -1653
rect 1477 -1653 1519 -1649
rect 1477 -1655 1490 -1653
rect 1411 -1670 1490 -1655
rect 1507 -1670 1519 -1653
rect 1536 -1659 1563 -1649
rect 1382 -1675 1519 -1670
rect 1443 -1686 1463 -1675
rect 1441 -1906 1461 -1895
rect 1380 -1911 1517 -1906
rect 1329 -1932 1363 -1922
rect 1380 -1928 1392 -1911
rect 1409 -1926 1488 -1911
rect 1409 -1928 1422 -1926
rect 1380 -1932 1422 -1928
rect 1475 -1928 1488 -1926
rect 1505 -1928 1517 -1911
rect 1475 -1932 1517 -1928
rect 1534 -1932 1561 -1922
rect 1329 -1951 1334 -1932
rect 1351 -1951 1363 -1932
rect 1534 -1951 1539 -1932
rect 1556 -1951 1561 -1932
rect 1329 -1961 1363 -1951
rect 1380 -1955 1422 -1951
rect 1380 -1972 1392 -1955
rect 1409 -1972 1422 -1955
rect 1380 -1977 1422 -1972
rect 1475 -1955 1517 -1951
rect 1475 -1972 1488 -1955
rect 1505 -1972 1517 -1955
rect 1534 -1961 1561 -1951
rect 1475 -1977 1517 -1972
rect 1390 -2004 1409 -1977
rect 1488 -2004 1507 -1977
rect 1380 -2009 1422 -2004
rect 1329 -2030 1363 -2020
rect 1380 -2026 1392 -2009
rect 1409 -2026 1422 -2009
rect 1380 -2030 1422 -2026
rect 1475 -2009 1517 -2004
rect 1475 -2026 1488 -2009
rect 1505 -2026 1517 -2009
rect 1475 -2030 1517 -2026
rect 1534 -2030 1561 -2020
rect 1329 -2049 1334 -2030
rect 1351 -2049 1363 -2030
rect 1534 -2049 1539 -2030
rect 1556 -2049 1561 -2030
rect 1329 -2059 1363 -2049
rect 1380 -2053 1422 -2049
rect 1380 -2070 1392 -2053
rect 1409 -2055 1422 -2053
rect 1475 -2053 1517 -2049
rect 1475 -2055 1488 -2053
rect 1409 -2070 1488 -2055
rect 1505 -2070 1517 -2053
rect 1534 -2059 1561 -2049
rect 1380 -2075 1517 -2070
rect 1441 -2086 1461 -2075
rect 1443 -2306 1463 -2295
rect 1382 -2311 1519 -2306
rect 1331 -2332 1365 -2322
rect 1382 -2328 1394 -2311
rect 1411 -2326 1490 -2311
rect 1411 -2328 1424 -2326
rect 1382 -2332 1424 -2328
rect 1477 -2328 1490 -2326
rect 1507 -2328 1519 -2311
rect 1477 -2332 1519 -2328
rect 1536 -2332 1563 -2322
rect 1331 -2351 1336 -2332
rect 1353 -2351 1365 -2332
rect 1536 -2351 1541 -2332
rect 1558 -2351 1563 -2332
rect 1331 -2361 1365 -2351
rect 1382 -2355 1424 -2351
rect 1382 -2372 1394 -2355
rect 1411 -2372 1424 -2355
rect 1382 -2377 1424 -2372
rect 1477 -2355 1519 -2351
rect 1477 -2372 1490 -2355
rect 1507 -2372 1519 -2355
rect 1536 -2361 1563 -2351
rect 1477 -2377 1519 -2372
rect 1392 -2404 1411 -2377
rect 1490 -2404 1509 -2377
rect 1382 -2409 1424 -2404
rect 1331 -2430 1365 -2420
rect 1382 -2426 1394 -2409
rect 1411 -2426 1424 -2409
rect 1382 -2430 1424 -2426
rect 1477 -2409 1519 -2404
rect 1477 -2426 1490 -2409
rect 1507 -2426 1519 -2409
rect 1477 -2430 1519 -2426
rect 1536 -2430 1563 -2420
rect 1331 -2449 1336 -2430
rect 1353 -2449 1365 -2430
rect 1536 -2449 1541 -2430
rect 1558 -2449 1563 -2430
rect 1331 -2459 1365 -2449
rect 1382 -2453 1424 -2449
rect 1382 -2470 1394 -2453
rect 1411 -2455 1424 -2453
rect 1477 -2453 1519 -2449
rect 1477 -2455 1490 -2453
rect 1411 -2470 1490 -2455
rect 1507 -2470 1519 -2453
rect 1536 -2459 1563 -2449
rect 1382 -2475 1519 -2470
rect 1443 -2486 1463 -2475
rect 1443 -2706 1463 -2695
rect 1382 -2711 1519 -2706
rect 1331 -2732 1365 -2722
rect 1382 -2728 1394 -2711
rect 1411 -2726 1490 -2711
rect 1411 -2728 1424 -2726
rect 1382 -2732 1424 -2728
rect 1477 -2728 1490 -2726
rect 1507 -2728 1519 -2711
rect 1477 -2732 1519 -2728
rect 1536 -2732 1563 -2722
rect 1331 -2751 1336 -2732
rect 1353 -2751 1365 -2732
rect 1536 -2751 1541 -2732
rect 1558 -2751 1563 -2732
rect 1331 -2761 1365 -2751
rect 1382 -2755 1424 -2751
rect 1382 -2772 1394 -2755
rect 1411 -2772 1424 -2755
rect 1382 -2777 1424 -2772
rect 1477 -2755 1519 -2751
rect 1477 -2772 1490 -2755
rect 1507 -2772 1519 -2755
rect 1536 -2761 1563 -2751
rect 1477 -2777 1519 -2772
rect 1392 -2804 1411 -2777
rect 1490 -2804 1509 -2777
rect 1382 -2809 1424 -2804
rect 1331 -2830 1365 -2820
rect 1382 -2826 1394 -2809
rect 1411 -2826 1424 -2809
rect 1382 -2830 1424 -2826
rect 1477 -2809 1519 -2804
rect 1477 -2826 1490 -2809
rect 1507 -2826 1519 -2809
rect 1477 -2830 1519 -2826
rect 1536 -2830 1563 -2820
rect 1331 -2849 1336 -2830
rect 1353 -2849 1365 -2830
rect 1536 -2849 1541 -2830
rect 1558 -2849 1563 -2830
rect 1331 -2859 1365 -2849
rect 1382 -2853 1424 -2849
rect 1382 -2870 1394 -2853
rect 1411 -2855 1424 -2853
rect 1477 -2853 1519 -2849
rect 1477 -2855 1490 -2853
rect 1411 -2870 1490 -2855
rect 1507 -2870 1519 -2853
rect 1536 -2859 1563 -2849
rect 1382 -2875 1519 -2870
rect 1443 -2886 1463 -2875
rect 1443 -3106 1463 -3095
rect 1382 -3111 1519 -3106
rect 1331 -3132 1365 -3122
rect 1382 -3128 1394 -3111
rect 1411 -3126 1490 -3111
rect 1411 -3128 1424 -3126
rect 1382 -3132 1424 -3128
rect 1477 -3128 1490 -3126
rect 1507 -3128 1519 -3111
rect 1477 -3132 1519 -3128
rect 1536 -3132 1563 -3122
rect 1331 -3151 1336 -3132
rect 1353 -3151 1365 -3132
rect 1536 -3151 1541 -3132
rect 1558 -3151 1563 -3132
rect 1331 -3161 1365 -3151
rect 1382 -3155 1424 -3151
rect 1382 -3172 1394 -3155
rect 1411 -3172 1424 -3155
rect 1382 -3177 1424 -3172
rect 1477 -3155 1519 -3151
rect 1477 -3172 1490 -3155
rect 1507 -3172 1519 -3155
rect 1536 -3161 1563 -3151
rect 1477 -3177 1519 -3172
rect 1392 -3204 1411 -3177
rect 1490 -3204 1509 -3177
rect 1382 -3209 1424 -3204
rect 1331 -3230 1365 -3220
rect 1382 -3226 1394 -3209
rect 1411 -3226 1424 -3209
rect 1382 -3230 1424 -3226
rect 1477 -3209 1519 -3204
rect 1477 -3226 1490 -3209
rect 1507 -3226 1519 -3209
rect 1477 -3230 1519 -3226
rect 1536 -3230 1563 -3220
rect 1331 -3249 1336 -3230
rect 1353 -3249 1365 -3230
rect 1536 -3249 1541 -3230
rect 1558 -3249 1563 -3230
rect 1331 -3259 1365 -3249
rect 1382 -3253 1424 -3249
rect 1382 -3270 1394 -3253
rect 1411 -3255 1424 -3253
rect 1477 -3253 1519 -3249
rect 1477 -3255 1490 -3253
rect 1411 -3270 1490 -3255
rect 1507 -3270 1519 -3253
rect 1536 -3259 1563 -3249
rect 1382 -3275 1519 -3270
rect 1443 -3286 1463 -3275
rect 1443 -3506 1463 -3495
rect 1382 -3511 1519 -3506
rect 1331 -3532 1365 -3522
rect 1382 -3528 1394 -3511
rect 1411 -3526 1490 -3511
rect 1411 -3528 1424 -3526
rect 1382 -3532 1424 -3528
rect 1477 -3528 1490 -3526
rect 1507 -3528 1519 -3511
rect 1477 -3532 1519 -3528
rect 1536 -3532 1563 -3522
rect 1331 -3551 1336 -3532
rect 1353 -3551 1365 -3532
rect 1536 -3551 1541 -3532
rect 1558 -3551 1563 -3532
rect 1331 -3561 1365 -3551
rect 1382 -3555 1424 -3551
rect 1382 -3572 1394 -3555
rect 1411 -3572 1424 -3555
rect 1382 -3577 1424 -3572
rect 1477 -3555 1519 -3551
rect 1477 -3572 1490 -3555
rect 1507 -3572 1519 -3555
rect 1536 -3561 1563 -3551
rect 1477 -3577 1519 -3572
rect 1392 -3604 1411 -3577
rect 1490 -3604 1509 -3577
rect 1382 -3609 1424 -3604
rect 1331 -3630 1365 -3620
rect 1382 -3626 1394 -3609
rect 1411 -3626 1424 -3609
rect 1382 -3630 1424 -3626
rect 1477 -3609 1519 -3604
rect 1477 -3626 1490 -3609
rect 1507 -3626 1519 -3609
rect 1477 -3630 1519 -3626
rect 1536 -3630 1563 -3620
rect 1331 -3649 1336 -3630
rect 1353 -3649 1365 -3630
rect 1536 -3649 1541 -3630
rect 1558 -3649 1563 -3630
rect 1331 -3659 1365 -3649
rect 1382 -3653 1424 -3649
rect 1382 -3670 1394 -3653
rect 1411 -3655 1424 -3653
rect 1477 -3653 1519 -3649
rect 1477 -3655 1490 -3653
rect 1411 -3670 1490 -3655
rect 1507 -3670 1519 -3653
rect 1536 -3659 1563 -3649
rect 1382 -3675 1519 -3670
rect 1443 -3686 1463 -3675
rect 23 -3798 87 -3771
rect 448 -3791 500 -3771
rect 135 -3797 155 -3791
rect 23 -3860 50 -3798
rect 131 -3837 155 -3797
rect 135 -3843 155 -3837
rect 448 -3853 477 -3791
rect 549 -3836 576 -3771
rect 869 -3798 935 -3770
rect 448 -3912 468 -3853
rect 869 -3865 896 -3798
rect 981 -3852 1001 -3782
<< viali >>
rect 1336 -351 1353 -332
rect 1541 -351 1558 -332
rect 1394 -372 1411 -355
rect 1490 -372 1507 -355
rect 1394 -426 1411 -409
rect 1490 -426 1507 -409
rect 1336 -449 1353 -430
rect 1541 -449 1558 -430
rect 1336 -751 1353 -732
rect 1541 -751 1558 -732
rect 1394 -772 1411 -755
rect 1490 -772 1507 -755
rect 1394 -826 1411 -809
rect 1490 -826 1507 -809
rect 1336 -849 1353 -830
rect 1541 -849 1558 -830
rect 1335 -1151 1352 -1132
rect 1540 -1151 1557 -1132
rect 1393 -1172 1410 -1155
rect 1489 -1172 1506 -1155
rect 1393 -1226 1410 -1209
rect 1489 -1226 1506 -1209
rect 1335 -1249 1352 -1230
rect 1540 -1249 1557 -1230
rect 1336 -1551 1353 -1532
rect 1541 -1551 1558 -1532
rect 1394 -1572 1411 -1555
rect 1490 -1572 1507 -1555
rect 1394 -1626 1411 -1609
rect 1490 -1626 1507 -1609
rect 1336 -1649 1353 -1630
rect 1541 -1649 1558 -1630
rect 1334 -1951 1351 -1932
rect 1539 -1951 1556 -1932
rect 1392 -1972 1409 -1955
rect 1488 -1972 1505 -1955
rect 1392 -2026 1409 -2009
rect 1488 -2026 1505 -2009
rect 1334 -2049 1351 -2030
rect 1539 -2049 1556 -2030
rect 1336 -2351 1353 -2332
rect 1541 -2351 1558 -2332
rect 1394 -2372 1411 -2355
rect 1490 -2372 1507 -2355
rect 1394 -2426 1411 -2409
rect 1490 -2426 1507 -2409
rect 1336 -2449 1353 -2430
rect 1541 -2449 1558 -2430
rect 1336 -2751 1353 -2732
rect 1541 -2751 1558 -2732
rect 1394 -2772 1411 -2755
rect 1490 -2772 1507 -2755
rect 1394 -2826 1411 -2809
rect 1490 -2826 1507 -2809
rect 1336 -2849 1353 -2830
rect 1541 -2849 1558 -2830
rect 1336 -3151 1353 -3132
rect 1541 -3151 1558 -3132
rect 1394 -3172 1411 -3155
rect 1490 -3172 1507 -3155
rect 1394 -3226 1411 -3209
rect 1490 -3226 1507 -3209
rect 1336 -3249 1353 -3230
rect 1541 -3249 1558 -3230
rect 1336 -3551 1353 -3532
rect 1541 -3551 1558 -3532
rect 1394 -3572 1411 -3555
rect 1490 -3572 1507 -3555
rect 1394 -3626 1411 -3609
rect 1490 -3626 1507 -3609
rect 1336 -3649 1353 -3630
rect 1541 -3649 1558 -3630
<< metal1 >>
rect 1250 153 1357 175
rect 1335 127 1357 153
rect 1252 107 1357 127
rect 1332 75 1357 107
rect 1335 61 1357 75
rect 1269 0 1425 23
rect 1383 -14 1425 0
rect 1332 -76 1354 -53
rect 1233 -96 1354 -76
rect 1332 -122 1354 -96
rect 1250 -144 1354 -122
rect 1272 -247 1356 -225
rect 1334 -273 1356 -247
rect 1272 -293 1356 -273
rect 1331 -322 1356 -293
rect 1331 -332 1359 -322
rect 1331 -351 1336 -332
rect 1353 -351 1359 -332
rect 1535 -332 1563 -322
rect 1331 -362 1359 -351
rect 1382 -355 1424 -349
rect 1382 -372 1394 -355
rect 1411 -372 1424 -355
rect 1382 -377 1424 -372
rect 1477 -355 1519 -348
rect 1477 -372 1490 -355
rect 1507 -372 1519 -355
rect 1535 -351 1541 -332
rect 1558 -351 1563 -332
rect 1535 -362 1563 -351
rect 1477 -377 1519 -372
rect 1272 -400 1424 -377
rect 1382 -409 1424 -400
rect 1331 -430 1359 -419
rect 1331 -449 1336 -430
rect 1353 -449 1359 -430
rect 1382 -426 1394 -409
rect 1411 -426 1424 -409
rect 1382 -432 1424 -426
rect 1477 -409 1519 -404
rect 1477 -426 1490 -409
rect 1507 -426 1519 -409
rect 1477 -433 1519 -426
rect 1535 -430 1563 -419
rect 1331 -459 1359 -449
rect 1535 -449 1541 -430
rect 1558 -449 1563 -430
rect 1535 -459 1563 -449
rect 1331 -476 1353 -459
rect 1272 -496 1353 -476
rect 1331 -522 1353 -496
rect 1272 -544 1353 -522
rect 1272 -647 1356 -625
rect 1334 -673 1356 -647
rect 1272 -693 1356 -673
rect 1331 -722 1356 -693
rect 1331 -732 1359 -722
rect 1331 -751 1336 -732
rect 1353 -751 1359 -732
rect 1535 -732 1563 -722
rect 1331 -762 1359 -751
rect 1382 -755 1424 -749
rect 1382 -772 1394 -755
rect 1411 -772 1424 -755
rect 1382 -777 1424 -772
rect 1477 -755 1519 -748
rect 1477 -772 1490 -755
rect 1507 -772 1519 -755
rect 1535 -751 1541 -732
rect 1558 -751 1563 -732
rect 1535 -762 1563 -751
rect 1477 -777 1519 -772
rect 1272 -800 1424 -777
rect 1382 -809 1424 -800
rect 1331 -830 1359 -819
rect 1331 -849 1336 -830
rect 1353 -849 1359 -830
rect 1382 -826 1394 -809
rect 1411 -826 1424 -809
rect 1382 -832 1424 -826
rect 1477 -809 1519 -804
rect 1477 -826 1490 -809
rect 1507 -826 1519 -809
rect 1477 -833 1519 -826
rect 1535 -830 1563 -819
rect 1331 -859 1359 -849
rect 1535 -849 1541 -830
rect 1558 -849 1563 -830
rect 1535 -859 1563 -849
rect 1331 -876 1353 -859
rect 1272 -896 1353 -876
rect 1331 -922 1353 -896
rect 1272 -944 1353 -922
rect 1271 -1047 1355 -1025
rect 1333 -1073 1355 -1047
rect 1271 -1093 1355 -1073
rect 1330 -1122 1355 -1093
rect 1330 -1132 1358 -1122
rect 1330 -1151 1335 -1132
rect 1352 -1151 1358 -1132
rect 1534 -1132 1562 -1122
rect 1330 -1162 1358 -1151
rect 1381 -1155 1423 -1149
rect 1381 -1172 1393 -1155
rect 1410 -1172 1423 -1155
rect 1381 -1177 1423 -1172
rect 1476 -1155 1518 -1148
rect 1476 -1172 1489 -1155
rect 1506 -1172 1518 -1155
rect 1534 -1151 1540 -1132
rect 1557 -1151 1562 -1132
rect 1534 -1162 1562 -1151
rect 1476 -1177 1518 -1172
rect 1271 -1200 1423 -1177
rect 1381 -1209 1423 -1200
rect 1330 -1230 1358 -1219
rect 1330 -1249 1335 -1230
rect 1352 -1249 1358 -1230
rect 1381 -1226 1393 -1209
rect 1410 -1226 1423 -1209
rect 1381 -1232 1423 -1226
rect 1476 -1209 1518 -1204
rect 1476 -1226 1489 -1209
rect 1506 -1226 1518 -1209
rect 1476 -1233 1518 -1226
rect 1534 -1230 1562 -1219
rect 1330 -1259 1358 -1249
rect 1534 -1249 1540 -1230
rect 1557 -1249 1562 -1230
rect 1534 -1259 1562 -1249
rect 1330 -1276 1352 -1259
rect 1271 -1296 1352 -1276
rect 1330 -1322 1352 -1296
rect 1271 -1344 1352 -1322
rect 1272 -1447 1356 -1425
rect 1334 -1473 1356 -1447
rect 1272 -1493 1356 -1473
rect 1331 -1522 1356 -1493
rect 1331 -1532 1359 -1522
rect 1331 -1551 1336 -1532
rect 1353 -1551 1359 -1532
rect 1535 -1532 1563 -1522
rect 1331 -1562 1359 -1551
rect 1382 -1555 1424 -1549
rect 1382 -1572 1394 -1555
rect 1411 -1572 1424 -1555
rect 1382 -1577 1424 -1572
rect 1477 -1555 1519 -1548
rect 1477 -1572 1490 -1555
rect 1507 -1572 1519 -1555
rect 1535 -1551 1541 -1532
rect 1558 -1551 1563 -1532
rect 1535 -1562 1563 -1551
rect 1477 -1577 1519 -1572
rect 1272 -1595 1424 -1577
rect 1089 -1600 1424 -1595
rect 1382 -1609 1424 -1600
rect 1331 -1630 1359 -1619
rect 1331 -1649 1336 -1630
rect 1353 -1649 1359 -1630
rect 1382 -1626 1394 -1609
rect 1411 -1626 1424 -1609
rect 1382 -1632 1424 -1626
rect 1477 -1609 1519 -1604
rect 1477 -1626 1490 -1609
rect 1507 -1626 1519 -1609
rect 1477 -1633 1519 -1626
rect 1535 -1630 1563 -1619
rect 1331 -1659 1359 -1649
rect 1535 -1649 1541 -1630
rect 1558 -1649 1563 -1630
rect 1535 -1659 1563 -1649
rect 1331 -1676 1353 -1659
rect 1272 -1696 1353 -1676
rect 1331 -1722 1353 -1696
rect 1272 -1744 1353 -1722
rect 1270 -1847 1354 -1825
rect 1332 -1873 1354 -1847
rect 1270 -1893 1354 -1873
rect 1329 -1922 1354 -1893
rect 1329 -1932 1357 -1922
rect 1329 -1951 1334 -1932
rect 1351 -1951 1357 -1932
rect 1533 -1932 1561 -1922
rect 1329 -1962 1357 -1951
rect 1380 -1955 1422 -1949
rect 1380 -1972 1392 -1955
rect 1409 -1972 1422 -1955
rect 1380 -1977 1422 -1972
rect 1475 -1955 1517 -1948
rect 1475 -1972 1488 -1955
rect 1505 -1972 1517 -1955
rect 1533 -1951 1539 -1932
rect 1556 -1951 1561 -1932
rect 1533 -1962 1561 -1951
rect 1475 -1977 1517 -1972
rect 1270 -1995 1422 -1977
rect 1089 -2000 1422 -1995
rect 1380 -2009 1422 -2000
rect 1329 -2030 1357 -2019
rect 1329 -2049 1334 -2030
rect 1351 -2049 1357 -2030
rect 1380 -2026 1392 -2009
rect 1409 -2026 1422 -2009
rect 1380 -2032 1422 -2026
rect 1475 -2009 1517 -2004
rect 1475 -2026 1488 -2009
rect 1505 -2026 1517 -2009
rect 1475 -2033 1517 -2026
rect 1533 -2030 1561 -2019
rect 1329 -2059 1357 -2049
rect 1533 -2049 1539 -2030
rect 1556 -2049 1561 -2030
rect 1533 -2059 1561 -2049
rect 1329 -2076 1351 -2059
rect 1270 -2096 1351 -2076
rect 1329 -2122 1351 -2096
rect 1270 -2144 1351 -2122
rect 1272 -2247 1356 -2225
rect 1334 -2273 1356 -2247
rect 1272 -2293 1356 -2273
rect 1331 -2322 1356 -2293
rect 1331 -2332 1359 -2322
rect 1331 -2351 1336 -2332
rect 1353 -2351 1359 -2332
rect 1535 -2332 1563 -2322
rect 1331 -2362 1359 -2351
rect 1382 -2355 1424 -2349
rect 1382 -2372 1394 -2355
rect 1411 -2372 1424 -2355
rect 1382 -2377 1424 -2372
rect 1477 -2355 1519 -2348
rect 1477 -2372 1490 -2355
rect 1507 -2372 1519 -2355
rect 1535 -2351 1541 -2332
rect 1558 -2351 1563 -2332
rect 1535 -2362 1563 -2351
rect 1477 -2377 1519 -2372
rect 1272 -2400 1424 -2377
rect 1382 -2409 1424 -2400
rect 1331 -2430 1359 -2419
rect 1331 -2449 1336 -2430
rect 1353 -2449 1359 -2430
rect 1382 -2426 1394 -2409
rect 1411 -2426 1424 -2409
rect 1382 -2432 1424 -2426
rect 1477 -2409 1519 -2404
rect 1477 -2426 1490 -2409
rect 1507 -2426 1519 -2409
rect 1477 -2433 1519 -2426
rect 1535 -2430 1563 -2419
rect 1331 -2459 1359 -2449
rect 1535 -2449 1541 -2430
rect 1558 -2449 1563 -2430
rect 1535 -2459 1563 -2449
rect 1331 -2476 1353 -2459
rect 1272 -2496 1353 -2476
rect 1331 -2522 1353 -2496
rect 1272 -2544 1353 -2522
rect 1272 -2647 1356 -2625
rect 1334 -2673 1356 -2647
rect 1272 -2693 1356 -2673
rect 1331 -2722 1356 -2693
rect 1331 -2732 1359 -2722
rect 1331 -2751 1336 -2732
rect 1353 -2751 1359 -2732
rect 1535 -2732 1563 -2722
rect 1331 -2762 1359 -2751
rect 1382 -2755 1424 -2749
rect 1382 -2772 1394 -2755
rect 1411 -2772 1424 -2755
rect 1382 -2777 1424 -2772
rect 1477 -2755 1519 -2748
rect 1477 -2772 1490 -2755
rect 1507 -2772 1519 -2755
rect 1535 -2751 1541 -2732
rect 1558 -2751 1563 -2732
rect 1535 -2762 1563 -2751
rect 1477 -2777 1519 -2772
rect 1272 -2800 1424 -2777
rect 1382 -2809 1424 -2800
rect 1331 -2830 1359 -2819
rect 1331 -2849 1336 -2830
rect 1353 -2849 1359 -2830
rect 1382 -2826 1394 -2809
rect 1411 -2826 1424 -2809
rect 1382 -2832 1424 -2826
rect 1477 -2809 1519 -2804
rect 1477 -2826 1490 -2809
rect 1507 -2826 1519 -2809
rect 1477 -2833 1519 -2826
rect 1535 -2830 1563 -2819
rect 1331 -2859 1359 -2849
rect 1535 -2849 1541 -2830
rect 1558 -2849 1563 -2830
rect 1535 -2859 1563 -2849
rect 1331 -2876 1353 -2859
rect 1272 -2896 1353 -2876
rect 1331 -2922 1353 -2896
rect 1272 -2944 1353 -2922
rect 1272 -3047 1356 -3025
rect 1334 -3073 1356 -3047
rect 1272 -3093 1356 -3073
rect 1331 -3122 1356 -3093
rect 1331 -3132 1359 -3122
rect 1331 -3151 1336 -3132
rect 1353 -3151 1359 -3132
rect 1535 -3132 1563 -3122
rect 1331 -3162 1359 -3151
rect 1382 -3155 1424 -3149
rect 1382 -3172 1394 -3155
rect 1411 -3172 1424 -3155
rect 1382 -3177 1424 -3172
rect 1477 -3155 1519 -3148
rect 1477 -3172 1490 -3155
rect 1507 -3172 1519 -3155
rect 1535 -3151 1541 -3132
rect 1558 -3151 1563 -3132
rect 1535 -3162 1563 -3151
rect 1477 -3177 1519 -3172
rect 1272 -3200 1424 -3177
rect 1382 -3209 1424 -3200
rect 1331 -3230 1359 -3219
rect 1331 -3249 1336 -3230
rect 1353 -3249 1359 -3230
rect 1382 -3226 1394 -3209
rect 1411 -3226 1424 -3209
rect 1382 -3232 1424 -3226
rect 1477 -3209 1519 -3204
rect 1477 -3226 1490 -3209
rect 1507 -3226 1519 -3209
rect 1477 -3233 1519 -3226
rect 1535 -3230 1563 -3219
rect 1331 -3259 1359 -3249
rect 1535 -3249 1541 -3230
rect 1558 -3249 1563 -3230
rect 1535 -3259 1563 -3249
rect 1331 -3276 1353 -3259
rect 1272 -3296 1353 -3276
rect 1331 -3322 1353 -3296
rect 1272 -3344 1353 -3322
rect 1272 -3447 1356 -3425
rect 1334 -3473 1356 -3447
rect 1272 -3493 1356 -3473
rect 1331 -3522 1356 -3493
rect 1331 -3532 1359 -3522
rect 1331 -3551 1336 -3532
rect 1353 -3551 1359 -3532
rect 1535 -3532 1563 -3522
rect 1331 -3562 1359 -3551
rect 1382 -3555 1424 -3549
rect 1382 -3572 1394 -3555
rect 1411 -3572 1424 -3555
rect 1382 -3577 1424 -3572
rect 1477 -3555 1519 -3548
rect 1477 -3572 1490 -3555
rect 1507 -3572 1519 -3555
rect 1535 -3551 1541 -3532
rect 1558 -3551 1563 -3532
rect 1535 -3562 1563 -3551
rect 1477 -3577 1519 -3572
rect 1272 -3600 1424 -3577
rect 1382 -3609 1424 -3600
rect 1331 -3630 1359 -3619
rect 1331 -3649 1336 -3630
rect 1353 -3649 1359 -3630
rect 1382 -3626 1394 -3609
rect 1411 -3626 1424 -3609
rect 1382 -3632 1424 -3626
rect 1477 -3609 1519 -3604
rect 1477 -3626 1490 -3609
rect 1507 -3626 1519 -3609
rect 1477 -3633 1519 -3626
rect 1535 -3630 1563 -3619
rect 1331 -3659 1359 -3649
rect 1535 -3649 1541 -3630
rect 1558 -3649 1563 -3630
rect 1535 -3659 1563 -3649
rect 1331 -3676 1353 -3659
rect 1272 -3696 1353 -3676
rect 1331 -3722 1353 -3696
rect 1272 -3744 1353 -3722
use buffer  buffer_0
timestamp 1640997824
transform 0 -1 255 1 0 -4088
box -14 -3 272 253
use buffer  buffer_1
timestamp 1640997824
transform 0 -1 679 1 0 -4088
box -14 -3 272 253
use buffer  buffer_2
timestamp 1640997824
transform 0 -1 1101 1 0 -4086
box -14 -3 272 253
use decoder_cell_0  decoder_cell_0_58
timestamp 1641069145
transform 1 0 1126 0 -1 -3416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_57
timestamp 1641069145
transform -1 0 994 0 -1 -3416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_62
timestamp 1641069145
transform 1 0 702 0 -1 -3416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_67
timestamp 1641069145
transform -1 0 146 0 -1 -3416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_66
array 0 1 212 0 0 229
timestamp 1641069145
transform 1 0 278 0 -1 -3416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_59
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 994 0 1 -3753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_63
timestamp 1641069145
transform 1 0 702 0 1 -3753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_64
timestamp 1641069145
transform -1 0 146 0 1 -3753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_65
array 0 1 212 0 0 229
timestamp 1641069145
transform 1 0 278 0 1 -3753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_54
timestamp 1641069145
transform 1 0 1126 0 1 -3353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_61
array 0 1 212 0 0 229
timestamp 1641069145
transform 1 0 278 0 1 -3353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_60
timestamp 1641069145
transform -1 0 146 0 1 -3353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_53
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 782 0 1 -3353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_50
timestamp 1641069145
transform 1 0 278 0 1 -2953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_49
timestamp 1641069145
transform -1 0 146 0 1 -2953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_43
array 0 3 -212 0 0 -229
timestamp 1641069145
transform -1 0 570 0 1 -2953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_52
timestamp 1641069145
transform -1 0 1206 0 -1 -3016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_51
timestamp 1641069145
transform 1 0 914 0 -1 -3016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_56
timestamp 1641069145
transform 1 0 278 0 -1 -3016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_55
timestamp 1641069145
transform -1 0 146 0 -1 -3016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_48
array 0 1 -212 0 0 229
timestamp 1641069145
transform -1 0 570 0 -1 -3016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_46
array 0 1 -212 0 0 229
timestamp 1641069145
transform -1 0 994 0 -1 -2616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_42
timestamp 1641069145
transform -1 0 570 0 -1 -2616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_47
timestamp 1641069145
transform 1 0 702 0 -1 -2616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_44
timestamp 1641069145
transform 1 0 278 0 -1 -2616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_45
timestamp 1641069145
transform -1 0 146 0 -1 -2616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_36
array 0 4 -212 0 0 229
timestamp 1641069145
transform -1 0 358 0 -1 -2216
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_37
timestamp 1641069145
transform -1 0 146 0 -1 -2216
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_41
timestamp 1641069145
transform -1 0 1206 0 1 -2553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_39
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 358 0 1 -2553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_40
array 0 1 212 0 0 -229
timestamp 1641069145
transform 1 0 702 0 1 -2553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_38
timestamp 1641069145
transform -1 0 146 0 1 -2553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_35
array 0 1 212 0 0 -229
timestamp 1641069145
transform 1 0 914 0 1 -2153
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_34
array 0 2 -212 0 0 -229
timestamp 1641069145
transform -1 0 358 0 1 -2153
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_32
timestamp 1641069145
transform -1 0 146 0 1 -2153
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_31
timestamp 1641069145
transform -1 0 146 0 -1 -1816
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_33
timestamp 1641069145
transform -1 0 358 0 -1 -1816
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_30
array 0 3 212 0 0 229
timestamp 1641069145
transform 1 0 490 0 -1 -1816
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_26
array 0 1 212 0 0 -229
timestamp 1641069145
transform 1 0 914 0 -1 -1416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_24
timestamp 1641069145
transform 1 0 66 0 -1 -1416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_25
array 0 2 -212 0 0 -229
timestamp 1641069145
transform -1 0 358 0 -1 -1416
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_27
timestamp 1641069145
transform 1 0 66 0 1 -1753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_29
array 0 3 212 0 0 229
timestamp 1641069145
transform 1 0 490 0 1 -1753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_28
timestamp 1641069145
transform -1 0 358 0 1 -1753
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_22
timestamp 1641069145
transform 1 0 66 0 1 -1353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_23
array 0 4 -212 0 0 229
timestamp 1641069145
transform -1 0 358 0 1 -1353
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_17
array 0 1 -212 0 0 229
timestamp 1641069145
transform -1 0 994 0 1 -953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_14
array 0 1 212 0 0 229
timestamp 1641069145
transform 1 0 66 0 1 -953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_16
timestamp 1641069145
transform 1 0 702 0 1 -953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_15
timestamp 1641069145
transform -1 0 570 0 1 -953
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_21
timestamp 1641069145
transform -1 0 1206 0 -1 -1016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_18
timestamp 1641069145
transform 1 0 66 0 -1 -1016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_19
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 358 0 -1 -1016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_20
array 0 1 212 0 0 -229
timestamp 1641069145
transform 1 0 702 0 -1 -1016
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_12
array 0 1 212 0 0 -229
timestamp 1641069145
transform 1 0 66 0 -1 -616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_13
array 0 3 -212 0 0 -229
timestamp 1641069145
transform -1 0 570 0 -1 -616
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_7
timestamp 1641069145
transform 1 0 1126 0 -1 -216
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_6
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 782 0 -1 -216
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_2
array 0 2 212 0 0 -229
timestamp 1641069145
transform 1 0 66 0 -1 -216
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_11
timestamp 1641069145
transform -1 0 1206 0 1 -553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_10
timestamp 1641069145
transform 1 0 914 0 1 -553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_9
array 0 1 -212 0 0 229
timestamp 1641069145
transform -1 0 570 0 1 -553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_8
array 0 1 212 0 0 229
timestamp 1641069145
transform 1 0 66 0 1 -553
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_5
timestamp 1641069145
transform 1 0 1126 0 1 -153
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_4
timestamp 1641069145
transform -1 0 994 0 1 -153
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_1
array 0 3 212 0 0 229
timestamp 1641069145
transform 1 0 66 0 1 -153
box -66 -45 146 184
use inv_lp  inv_lp_1
timestamp 1640995782
transform 0 -1 1522 -1 0 -43
box -61 -42 50 190
use decoder_cell_0  decoder_cell_0_3
array 0 1 -212 0 0 -229
timestamp 1641069145
transform -1 0 994 0 -1 184
box -66 -45 146 184
use decoder_cell_0  decoder_cell_0_0
array 0 3 212 0 0 -229
timestamp 1641069145
transform 1 0 66 0 -1 184
box -66 -45 146 184
use inv_lp  inv_lp_0
timestamp 1640995782
transform 0 -1 1522 1 0 62
box -61 -42 50 190
use buffer  buffer_3
timestamp 1640997824
transform 0 -1 466 -1 0 526
box -14 -3 272 253
use buffer  buffer_4
timestamp 1640997824
transform 0 -1 890 -1 0 525
box -14 -3 272 253
use buffer  buffer_5
timestamp 1640997824
transform 0 -1 1312 -1 0 526
box -14 -3 272 253
<< end >>
