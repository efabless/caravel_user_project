VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_2kbyte_1rw1r_32x512_8
   CLASS BLOCK ;
   SIZE 679.02 BY 413.14 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.56 0.0 113.94 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.0 0.0 119.38 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.12 0.0 125.5 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 0.0 130.94 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.0 0.0 136.38 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.36 0.0 154.74 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 0.0 160.18 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.24 0.0 165.62 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.48 0.0 177.86 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.92 0.0 183.3 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.36 0.0 188.74 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 0.0 195.54 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.72 0.0 207.1 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.16 0.0 212.54 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.84 0.0 247.22 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 0.0 259.46 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.52 0.0 264.9 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 0.0 270.34 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 0.0 277.14 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.88 0.0 283.26 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.76 0.0 294.14 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.2 0.0 78.58 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.64 0.0 84.02 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 139.4 0.38 139.78 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.24 0.38 148.62 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.36 0.38 154.74 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 162.52 0.38 162.9 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.96 0.38 168.34 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 177.48 0.38 177.86 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 182.92 0.38 183.3 ;
      END
   END addr0[8]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  596.36 412.76 596.74 413.14 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  590.24 412.76 590.62 413.14 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 95.2 679.02 95.58 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 87.04 679.02 87.42 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 80.24 679.02 80.62 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 72.76 679.02 73.14 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 66.64 679.02 67.02 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  614.04 0.0 614.42 0.38 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  614.72 0.0 615.1 0.38 ;
      END
   END addr1[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 38.76 0.38 39.14 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  678.64 394.4 679.02 394.78 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 48.28 0.38 48.66 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 0.38 40.5 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  652.12 412.76 652.5 413.14 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.08 0.0 89.46 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.88 0.0 96.26 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  100.64 0.0 101.02 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.76 0.0 107.14 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 0.0 152.02 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 0.0 166.3 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 0.0 178.54 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 0.0 190.78 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.96 0.0 253.34 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 0.0 290.74 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  315.52 0.0 315.9 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 0.0 328.14 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  339.32 0.0 339.7 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  352.92 0.0 353.3 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.16 0.0 365.54 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 0.0 377.78 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  390.32 0.0 390.7 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  402.56 0.0 402.94 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 0.0 415.86 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  427.72 0.0 428.1 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  440.64 0.0 441.02 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 0.0 453.26 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  465.12 0.0 465.5 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  477.36 0.0 477.74 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.28 0.0 490.66 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  502.52 0.0 502.9 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  514.76 0.0 515.14 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  527.68 0.0 528.06 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 412.76 141.82 413.14 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.0 412.76 153.38 413.14 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.24 412.76 165.62 413.14 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 412.76 179.22 413.14 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.4 412.76 190.78 413.14 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 412.76 203.7 413.14 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 412.76 215.94 413.14 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 412.76 228.86 413.14 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.72 412.76 241.1 413.14 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 412.76 254.02 413.14 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 412.76 266.26 413.14 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 412.76 279.18 413.14 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.36 412.76 290.74 413.14 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 412.76 302.98 413.14 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 412.76 316.58 413.14 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.44 412.76 328.82 413.14 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.68 412.76 341.06 413.14 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  352.92 412.76 353.3 413.14 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.84 412.76 366.22 413.14 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 412.76 377.78 413.14 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.0 412.76 391.38 413.14 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  403.24 412.76 403.62 413.14 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 412.76 415.86 413.14 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  427.72 412.76 428.1 413.14 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  439.96 412.76 440.34 413.14 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 412.76 453.26 413.14 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  465.8 412.76 466.18 413.14 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  478.04 412.76 478.42 413.14 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.28 412.76 490.66 413.14 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  503.2 412.76 503.58 413.14 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  514.76 412.76 515.14 413.14 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  528.36 412.76 528.74 413.14 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  1.36 1.36 677.66 3.1 ;
         LAYER met4 ;
         RECT  675.92 1.36 677.66 411.78 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 411.78 ;
         LAYER met3 ;
         RECT  1.36 410.04 677.66 411.78 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 674.26 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 408.38 ;
         LAYER met3 ;
         RECT  4.76 406.64 674.26 408.38 ;
         LAYER met4 ;
         RECT  672.52 4.76 674.26 408.38 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 678.4 412.52 ;
   LAYER  met2 ;
      RECT  0.62 0.62 678.4 412.52 ;
   LAYER  met3 ;
      RECT  0.98 138.8 678.4 140.38 ;
      RECT  0.62 140.38 0.98 147.64 ;
      RECT  0.62 149.22 0.98 153.76 ;
      RECT  0.62 155.34 0.98 161.92 ;
      RECT  0.62 163.5 0.98 167.36 ;
      RECT  0.62 168.94 0.98 176.88 ;
      RECT  0.62 178.46 0.98 182.32 ;
      RECT  0.98 94.6 678.04 96.18 ;
      RECT  0.98 96.18 678.04 138.8 ;
      RECT  678.04 96.18 678.4 138.8 ;
      RECT  678.04 88.02 678.4 94.6 ;
      RECT  678.04 81.22 678.4 86.44 ;
      RECT  678.04 73.74 678.4 79.64 ;
      RECT  678.04 67.62 678.4 72.16 ;
      RECT  0.98 140.38 678.04 393.8 ;
      RECT  0.98 393.8 678.04 395.38 ;
      RECT  678.04 140.38 678.4 393.8 ;
      RECT  0.62 49.26 0.98 138.8 ;
      RECT  0.62 41.1 0.98 47.68 ;
      RECT  0.98 0.62 678.04 0.76 ;
      RECT  678.04 0.62 678.26 0.76 ;
      RECT  678.04 3.7 678.26 66.04 ;
      RECT  678.26 0.62 678.4 0.76 ;
      RECT  678.26 0.76 678.4 3.7 ;
      RECT  678.26 3.7 678.4 66.04 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 38.16 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 38.16 ;
      RECT  0.62 183.9 0.76 409.44 ;
      RECT  0.62 409.44 0.76 412.38 ;
      RECT  0.62 412.38 0.76 412.52 ;
      RECT  0.76 183.9 0.98 409.44 ;
      RECT  0.76 412.38 0.98 412.52 ;
      RECT  0.98 412.38 678.04 412.52 ;
      RECT  678.04 395.38 678.26 409.44 ;
      RECT  678.04 412.38 678.26 412.52 ;
      RECT  678.26 395.38 678.4 409.44 ;
      RECT  678.26 409.44 678.4 412.38 ;
      RECT  678.26 412.38 678.4 412.52 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 94.6 ;
      RECT  4.16 3.7 674.86 4.16 ;
      RECT  4.16 7.1 674.86 94.6 ;
      RECT  674.86 3.7 678.04 4.16 ;
      RECT  674.86 4.16 678.04 7.1 ;
      RECT  674.86 7.1 678.04 94.6 ;
      RECT  0.98 395.38 4.16 406.04 ;
      RECT  0.98 406.04 4.16 408.98 ;
      RECT  0.98 408.98 4.16 409.44 ;
      RECT  4.16 395.38 674.86 406.04 ;
      RECT  4.16 408.98 674.86 409.44 ;
      RECT  674.86 395.38 678.04 406.04 ;
      RECT  674.86 406.04 678.04 408.98 ;
      RECT  674.86 408.98 678.04 409.44 ;
   LAYER  met4 ;
      RECT  112.96 0.98 114.54 412.52 ;
      RECT  114.54 0.62 118.4 0.98 ;
      RECT  119.98 0.62 124.52 0.98 ;
      RECT  126.1 0.62 129.96 0.98 ;
      RECT  131.54 0.62 135.4 0.98 ;
      RECT  142.42 0.62 147.64 0.98 ;
      RECT  155.34 0.62 159.2 0.98 ;
      RECT  160.78 0.62 164.64 0.98 ;
      RECT  171.66 0.62 176.88 0.98 ;
      RECT  183.9 0.62 187.76 0.98 ;
      RECT  196.14 0.62 200.68 0.98 ;
      RECT  207.7 0.62 211.56 0.98 ;
      RECT  218.58 0.62 223.8 0.98 ;
      RECT  230.82 0.62 235.36 0.98 ;
      RECT  242.38 0.62 246.24 0.98 ;
      RECT  254.62 0.62 258.48 0.98 ;
      RECT  260.06 0.62 263.92 0.98 ;
      RECT  270.94 0.62 276.16 0.98 ;
      RECT  283.86 0.62 287.72 0.98 ;
      RECT  79.18 0.62 83.04 0.98 ;
      RECT  114.54 0.98 595.76 412.16 ;
      RECT  595.76 0.98 597.34 412.16 ;
      RECT  591.22 412.16 595.76 412.52 ;
      RECT  597.34 412.16 651.52 412.52 ;
      RECT  84.62 0.62 88.48 0.98 ;
      RECT  90.06 0.62 95.28 0.98 ;
      RECT  96.86 0.62 100.04 0.98 ;
      RECT  101.62 0.62 106.16 0.98 ;
      RECT  107.74 0.62 112.96 0.98 ;
      RECT  136.98 0.62 138.8 0.98 ;
      RECT  140.38 0.62 140.84 0.98 ;
      RECT  149.22 0.62 151.04 0.98 ;
      RECT  152.62 0.62 153.76 0.98 ;
      RECT  166.9 0.62 170.08 0.98 ;
      RECT  179.14 0.62 182.32 0.98 ;
      RECT  189.34 0.62 189.8 0.98 ;
      RECT  191.38 0.62 194.56 0.98 ;
      RECT  202.26 0.62 202.72 0.98 ;
      RECT  204.3 0.62 206.12 0.98 ;
      RECT  213.14 0.62 214.96 0.98 ;
      RECT  216.54 0.62 217.0 0.98 ;
      RECT  225.38 0.62 227.2 0.98 ;
      RECT  228.78 0.62 229.24 0.98 ;
      RECT  236.94 0.62 238.76 0.98 ;
      RECT  240.34 0.62 240.8 0.98 ;
      RECT  247.82 0.62 252.36 0.98 ;
      RECT  266.86 0.62 269.36 0.98 ;
      RECT  279.1 0.62 282.28 0.98 ;
      RECT  289.3 0.62 289.76 0.98 ;
      RECT  291.34 0.62 293.16 0.98 ;
      RECT  294.74 0.62 302.0 0.98 ;
      RECT  303.58 0.62 314.92 0.98 ;
      RECT  316.5 0.62 327.16 0.98 ;
      RECT  328.74 0.62 338.72 0.98 ;
      RECT  340.3 0.62 352.32 0.98 ;
      RECT  353.9 0.62 364.56 0.98 ;
      RECT  366.14 0.62 376.8 0.98 ;
      RECT  378.38 0.62 389.72 0.98 ;
      RECT  391.3 0.62 401.96 0.98 ;
      RECT  403.54 0.62 414.88 0.98 ;
      RECT  416.46 0.62 427.12 0.98 ;
      RECT  428.7 0.62 440.04 0.98 ;
      RECT  441.62 0.62 452.28 0.98 ;
      RECT  453.86 0.62 464.52 0.98 ;
      RECT  466.1 0.62 476.76 0.98 ;
      RECT  478.34 0.62 489.68 0.98 ;
      RECT  491.26 0.62 501.92 0.98 ;
      RECT  503.5 0.62 514.16 0.98 ;
      RECT  515.74 0.62 527.08 0.98 ;
      RECT  528.66 0.62 613.44 0.98 ;
      RECT  114.54 412.16 140.84 412.52 ;
      RECT  142.42 412.16 152.4 412.52 ;
      RECT  153.98 412.16 164.64 412.52 ;
      RECT  166.22 412.16 178.24 412.52 ;
      RECT  179.82 412.16 189.8 412.52 ;
      RECT  191.38 412.16 202.72 412.52 ;
      RECT  204.3 412.16 214.96 412.52 ;
      RECT  216.54 412.16 227.88 412.52 ;
      RECT  229.46 412.16 240.12 412.52 ;
      RECT  241.7 412.16 253.04 412.52 ;
      RECT  254.62 412.16 265.28 412.52 ;
      RECT  266.86 412.16 278.2 412.52 ;
      RECT  279.78 412.16 289.76 412.52 ;
      RECT  291.34 412.16 302.0 412.52 ;
      RECT  303.58 412.16 315.6 412.52 ;
      RECT  317.18 412.16 327.84 412.52 ;
      RECT  329.42 412.16 340.08 412.52 ;
      RECT  341.66 412.16 352.32 412.52 ;
      RECT  353.9 412.16 365.24 412.52 ;
      RECT  366.82 412.16 376.8 412.52 ;
      RECT  378.38 412.16 390.4 412.52 ;
      RECT  391.98 412.16 402.64 412.52 ;
      RECT  404.22 412.16 414.88 412.52 ;
      RECT  416.46 412.16 427.12 412.52 ;
      RECT  428.7 412.16 439.36 412.52 ;
      RECT  440.94 412.16 452.28 412.52 ;
      RECT  453.86 412.16 465.2 412.52 ;
      RECT  466.78 412.16 477.44 412.52 ;
      RECT  479.02 412.16 489.68 412.52 ;
      RECT  491.26 412.16 502.6 412.52 ;
      RECT  504.18 412.16 514.16 412.52 ;
      RECT  515.74 412.16 527.76 412.52 ;
      RECT  529.34 412.16 589.64 412.52 ;
      RECT  678.26 0.98 678.4 412.16 ;
      RECT  615.7 0.62 675.32 0.76 ;
      RECT  615.7 0.76 675.32 0.98 ;
      RECT  675.32 0.62 678.26 0.76 ;
      RECT  678.26 0.62 678.4 0.76 ;
      RECT  678.26 0.76 678.4 0.98 ;
      RECT  653.1 412.16 675.32 412.38 ;
      RECT  653.1 412.38 675.32 412.52 ;
      RECT  675.32 412.38 678.26 412.52 ;
      RECT  678.26 412.16 678.4 412.38 ;
      RECT  678.26 412.38 678.4 412.52 ;
      RECT  0.62 0.98 0.76 412.38 ;
      RECT  0.62 412.38 0.76 412.52 ;
      RECT  0.76 412.38 3.7 412.52 ;
      RECT  3.7 412.38 112.96 412.52 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 77.6 0.76 ;
      RECT  3.7 0.76 77.6 0.98 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 408.98 ;
      RECT  3.7 408.98 4.16 412.38 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 408.98 7.1 412.38 ;
      RECT  7.1 0.98 112.96 4.16 ;
      RECT  7.1 4.16 112.96 408.98 ;
      RECT  7.1 408.98 112.96 412.38 ;
      RECT  597.34 0.98 671.92 4.16 ;
      RECT  597.34 4.16 671.92 408.98 ;
      RECT  597.34 408.98 671.92 412.16 ;
      RECT  671.92 0.98 674.86 4.16 ;
      RECT  671.92 408.98 674.86 412.16 ;
      RECT  674.86 0.98 675.32 4.16 ;
      RECT  674.86 4.16 675.32 408.98 ;
      RECT  674.86 408.98 675.32 412.16 ;
   END
END    sky130_sram_2kbyte_1rw1r_32x512_8
END    LIBRARY
