magic
tech sky130A
timestamp 1641059315
<< nwell >>
rect -158 421 -3 526
rect -158 379 -72 421
<< nmos >>
rect -140 233 60 248
rect -140 126 60 141
rect -140 21 60 36
rect -140 -86 60 -71
rect -140 -195 60 -180
rect -140 -302 60 -287
rect -140 -407 60 -392
rect -140 -514 60 -499
rect -140 -616 60 -601
rect -140 -721 60 -706
rect -140 -828 60 -813
<< pmos >>
rect -140 436 -90 451
<< ndiff >>
rect -140 330 60 343
rect -140 259 -131 330
rect 48 259 60 330
rect -140 248 60 259
rect -140 222 60 233
rect -140 151 -129 222
rect 50 151 60 222
rect -140 141 60 151
rect -140 116 60 126
rect -140 45 -129 116
rect 50 45 60 116
rect -140 36 60 45
rect -140 8 60 21
rect -140 -63 -129 8
rect 50 -63 60 8
rect -140 -71 60 -63
rect -140 -99 60 -86
rect -140 -170 -129 -99
rect 50 -170 60 -99
rect -140 -180 60 -170
rect -140 -204 60 -195
rect -140 -275 -129 -204
rect 50 -275 60 -204
rect -140 -287 60 -275
rect -140 -311 60 -302
rect -140 -382 -130 -311
rect 49 -382 60 -311
rect -140 -392 60 -382
rect -140 -418 60 -407
rect -140 -489 -129 -418
rect 50 -489 60 -418
rect -140 -499 60 -489
rect -140 -523 60 -514
rect -140 -592 -130 -523
rect 49 -592 60 -523
rect -140 -601 60 -592
rect -140 -624 60 -616
rect -140 -700 -130 -624
rect 49 -700 60 -624
rect -140 -706 60 -700
rect -140 -728 60 -721
rect -140 -804 -130 -728
rect 49 -804 60 -728
rect -140 -813 60 -804
rect -140 -838 60 -828
rect -140 -914 -129 -838
rect 50 -914 60 -838
rect -140 -923 60 -914
<< pdiff >>
rect -140 481 -90 490
rect -140 464 -126 481
rect -100 464 -90 481
rect -140 451 -90 464
rect -140 424 -90 436
rect -140 407 -126 424
rect -100 407 -90 424
rect -140 397 -90 407
<< ndiffc >>
rect -131 259 48 330
rect -129 151 50 222
rect -129 45 50 116
rect -129 -63 50 8
rect -129 -170 50 -99
rect -129 -275 50 -204
rect -130 -382 49 -311
rect -129 -489 50 -418
rect -130 -592 49 -523
rect -130 -700 49 -624
rect -130 -804 49 -728
rect -129 -914 50 -838
<< pdiffc >>
rect -126 464 -100 481
rect -126 407 -100 424
<< psubdiff >>
rect -412 384 -321 412
rect -412 345 -387 384
rect -352 345 -321 384
rect -412 317 -321 345
<< nsubdiff >>
rect -62 488 -21 500
rect -62 471 -49 488
rect -32 471 -21 488
rect -62 458 -21 471
<< psubdiffcont >>
rect -387 345 -352 384
<< nsubdiffcont >>
rect -49 471 -32 488
<< poly >>
rect -193 451 -156 460
rect -193 434 -184 451
rect -165 436 -140 451
rect -90 436 -65 451
rect -165 434 -156 436
rect -193 425 -156 434
rect -193 249 -158 257
rect -193 232 -185 249
rect -166 248 -158 249
rect -166 233 -140 248
rect 60 233 85 248
rect -166 232 -158 233
rect -193 224 -158 232
rect -193 141 -158 149
rect -193 124 -186 141
rect -167 126 -140 141
rect 60 126 85 141
rect -167 124 -158 126
rect -193 116 -158 124
rect -193 37 -158 45
rect -193 20 -184 37
rect -165 36 -158 37
rect -165 21 -140 36
rect 60 21 85 36
rect -165 20 -158 21
rect -193 12 -158 20
rect -193 -70 -158 -62
rect -193 -87 -184 -70
rect -165 -71 -158 -70
rect -165 -86 -140 -71
rect 60 -86 85 -71
rect -165 -87 -158 -86
rect -193 -95 -158 -87
rect -193 -180 -158 -172
rect -193 -197 -185 -180
rect -166 -195 -140 -180
rect 60 -195 85 -180
rect -166 -197 -158 -195
rect -193 -205 -158 -197
rect -193 -286 -158 -278
rect -193 -303 -185 -286
rect -166 -287 -158 -286
rect -166 -302 -140 -287
rect 60 -302 85 -287
rect -166 -303 -158 -302
rect -193 -311 -158 -303
rect -193 -391 -158 -383
rect -193 -408 -185 -391
rect -166 -392 -158 -391
rect -166 -407 -140 -392
rect 60 -407 85 -392
rect -166 -408 -158 -407
rect -193 -416 -158 -408
rect -193 -498 -158 -490
rect -193 -515 -186 -498
rect -167 -499 -158 -498
rect -167 -514 -140 -499
rect 60 -514 85 -499
rect -167 -515 -158 -514
rect -193 -523 -158 -515
rect -193 -600 -158 -592
rect -193 -617 -185 -600
rect -166 -601 -158 -600
rect -166 -616 -140 -601
rect 60 -616 85 -601
rect -166 -617 -158 -616
rect -193 -625 -158 -617
rect -193 -704 -158 -696
rect -193 -721 -185 -704
rect -166 -706 -158 -704
rect -166 -721 -140 -706
rect 60 -721 85 -706
rect -193 -729 -158 -721
rect -193 -812 -158 -804
rect -193 -829 -185 -812
rect -166 -813 -158 -812
rect -166 -828 -140 -813
rect 60 -828 85 -813
rect -166 -829 -158 -828
rect -193 -837 -158 -829
<< polycont >>
rect -184 434 -165 451
rect -185 232 -166 249
rect -186 124 -167 141
rect -184 20 -165 37
rect -184 -87 -165 -70
rect -185 -197 -166 -180
rect -185 -303 -166 -286
rect -185 -408 -166 -391
rect -186 -515 -167 -498
rect -185 -617 -166 -600
rect -185 -721 -166 -704
rect -185 -829 -166 -812
<< locali >>
rect -138 489 -90 490
rect -62 489 -21 500
rect -138 488 -21 489
rect -138 481 -49 488
rect -138 464 -126 481
rect -100 471 -49 481
rect -32 471 -21 488
rect -100 464 -21 471
rect -138 461 -21 464
rect -256 451 -156 460
rect -138 455 -90 461
rect -62 458 -21 461
rect -256 434 -184 451
rect -165 434 -156 451
rect -256 425 -156 434
rect -138 431 -90 432
rect -256 424 -192 425
rect -138 424 171 431
rect -412 384 -321 412
rect -412 345 -387 384
rect -352 374 -321 384
rect -256 374 -220 424
rect -138 407 -126 424
rect -100 407 171 424
rect -138 398 171 407
rect -138 397 -90 398
rect -352 347 -220 374
rect -352 345 -321 347
rect -412 317 -321 345
rect -256 202 -220 347
rect -138 330 60 343
rect -138 259 -131 330
rect 48 309 60 330
rect 100 309 142 398
rect 48 267 142 309
rect 48 259 60 267
rect -193 249 -158 257
rect -138 250 60 259
rect -193 232 -185 249
rect -166 232 -158 249
rect -193 224 -158 232
rect -137 222 60 231
rect -137 202 -129 222
rect -256 166 -129 202
rect -256 -7 -220 166
rect -141 165 -129 166
rect -137 151 -129 165
rect 50 151 60 222
rect -193 141 -158 149
rect -137 143 60 151
rect -193 124 -186 141
rect -167 124 -158 141
rect -193 116 -158 124
rect -138 116 60 124
rect -138 45 -129 116
rect 50 109 60 116
rect 100 109 142 267
rect 50 67 142 109
rect 50 45 60 67
rect -193 37 -158 45
rect -138 38 60 45
rect -193 20 -184 37
rect -165 20 -158 37
rect -193 12 -158 20
rect -138 8 60 19
rect -138 -7 -129 8
rect -256 -43 -129 -7
rect -256 -224 -220 -43
rect -193 -70 -158 -62
rect -138 -63 -129 -43
rect 50 -63 60 8
rect -138 -69 60 -63
rect -193 -87 -184 -70
rect -165 -87 -158 -70
rect -193 -95 -158 -87
rect -138 -99 60 -88
rect -138 -170 -129 -99
rect 50 -114 60 -99
rect 100 -114 142 67
rect 50 -156 142 -114
rect 50 -170 60 -156
rect -193 -180 -158 -172
rect -138 -178 60 -170
rect -193 -197 -185 -180
rect -166 -197 -158 -180
rect -193 -205 -158 -197
rect -138 -204 60 -197
rect -138 -224 -129 -204
rect -256 -260 -129 -224
rect -256 -435 -220 -260
rect -138 -275 -129 -260
rect 50 -275 60 -204
rect -193 -286 -158 -278
rect -138 -285 60 -275
rect -193 -303 -185 -286
rect -166 -303 -158 -286
rect -193 -311 -158 -303
rect -138 -311 60 -304
rect -138 -382 -130 -311
rect 49 -339 60 -311
rect 100 -339 142 -156
rect 49 -381 142 -339
rect 49 -382 60 -381
rect -193 -391 -158 -383
rect -138 -390 60 -382
rect -193 -408 -185 -391
rect -166 -408 -158 -391
rect -193 -416 -158 -408
rect -138 -418 60 -409
rect -138 -435 -129 -418
rect -256 -471 -129 -435
rect -256 -644 -220 -471
rect -138 -489 -129 -471
rect 50 -489 60 -418
rect -193 -498 -158 -490
rect -138 -497 60 -489
rect -193 -515 -186 -498
rect -167 -515 -158 -498
rect -193 -523 -158 -515
rect -138 -523 60 -516
rect -138 -592 -130 -523
rect 49 -535 60 -523
rect 100 -535 142 -381
rect 49 -577 142 -535
rect 49 -592 60 -577
rect -193 -600 -158 -592
rect -138 -599 60 -592
rect -193 -617 -185 -600
rect -166 -617 -158 -600
rect -193 -625 -158 -617
rect -138 -624 60 -618
rect -138 -644 -130 -624
rect -256 -678 -130 -644
rect -256 -859 -220 -678
rect -140 -680 -130 -678
rect -193 -704 -158 -696
rect -138 -700 -130 -680
rect 49 -700 60 -624
rect -138 -704 60 -700
rect -193 -721 -185 -704
rect -166 -721 -158 -704
rect -193 -729 -158 -721
rect -138 -728 60 -723
rect -138 -804 -130 -728
rect 49 -744 60 -728
rect 100 -744 142 -577
rect 49 -804 142 -744
rect -193 -812 -158 -804
rect -138 -805 142 -804
rect -138 -811 60 -805
rect -193 -829 -185 -812
rect -166 -829 -158 -812
rect -193 -837 -158 -829
rect -138 -838 60 -830
rect -138 -859 -129 -838
rect -256 -914 -129 -859
rect 50 -914 60 -838
rect -256 -920 60 -914
rect -138 -921 60 -920
<< viali >>
rect -126 464 -100 481
rect -184 434 -165 451
rect -80 280 -12 311
rect -185 232 -166 249
rect -75 172 -7 203
rect -186 124 -167 141
rect -77 65 -9 96
rect -184 20 -165 37
rect -77 -45 -9 -14
rect -184 -87 -165 -70
rect -74 -151 -6 -120
rect -185 -197 -166 -180
rect -78 -254 -10 -223
rect -185 -303 -166 -286
rect -70 -361 -2 -330
rect -185 -408 -166 -391
rect -74 -468 -5 -440
rect -186 -515 -167 -498
rect -80 -573 -12 -545
rect -185 -617 -166 -600
rect -83 -679 0 -646
rect -185 -721 -166 -704
rect -79 -783 -6 -752
rect -185 -829 -166 -812
rect -76 -891 -4 -860
<< metal1 >>
rect -134 490 -107 518
rect -138 481 -90 490
rect -138 464 -126 481
rect -100 464 -90 481
rect -193 460 -156 461
rect -261 451 -156 460
rect -138 455 -90 464
rect -261 434 -184 451
rect -165 434 -156 451
rect -261 425 -156 434
rect -261 424 -157 425
rect -138 311 60 343
rect -138 280 -80 311
rect -12 280 60 311
rect -261 249 -158 257
rect -138 250 60 280
rect -261 232 -185 249
rect -166 232 -158 249
rect -261 224 -158 232
rect -137 203 60 231
rect -137 172 -75 203
rect -7 172 60 203
rect -260 141 -158 149
rect -137 143 60 172
rect -260 124 -186 141
rect -167 124 -158 141
rect -260 116 -158 124
rect -260 115 -161 116
rect -138 96 60 124
rect -138 65 -77 96
rect -9 65 60 96
rect -261 45 -163 46
rect -261 37 -158 45
rect -138 38 60 65
rect -261 20 -184 37
rect -165 20 -158 37
rect -261 12 -158 20
rect -138 -14 60 19
rect -138 -45 -77 -14
rect -9 -45 60 -14
rect -261 -62 -169 -61
rect -261 -70 -158 -62
rect -138 -69 60 -45
rect -261 -87 -184 -70
rect -165 -87 -158 -70
rect -261 -95 -158 -87
rect -138 -120 60 -88
rect -138 -151 -74 -120
rect -6 -151 60 -120
rect -261 -180 -158 -172
rect -138 -178 60 -151
rect -261 -197 -185 -180
rect -166 -197 -158 -180
rect -261 -205 -158 -197
rect -261 -206 -165 -205
rect -137 -223 60 -197
rect -137 -254 -78 -223
rect -10 -254 60 -223
rect -261 -278 -168 -277
rect -261 -286 -158 -278
rect -137 -285 60 -254
rect -261 -303 -185 -286
rect -166 -303 -158 -286
rect -261 -311 -158 -303
rect -138 -330 60 -305
rect -138 -361 -70 -330
rect -2 -361 60 -330
rect -261 -391 -158 -383
rect -138 -391 60 -361
rect -261 -408 -185 -391
rect -166 -408 -158 -391
rect -261 -416 -158 -408
rect -261 -417 -166 -416
rect -138 -440 60 -410
rect -138 -468 -74 -440
rect -5 -468 60 -440
rect -261 -498 -158 -490
rect -138 -496 60 -468
rect -261 -515 -186 -498
rect -167 -515 -158 -498
rect -261 -523 -158 -515
rect -261 -524 -167 -523
rect -138 -545 60 -516
rect -138 -573 -80 -545
rect -12 -573 60 -545
rect -261 -592 -163 -591
rect -261 -600 -158 -592
rect -138 -598 60 -573
rect -261 -617 -185 -600
rect -166 -617 -158 -600
rect -261 -625 -158 -617
rect -138 -646 61 -618
rect -138 -679 -83 -646
rect 0 -679 61 -646
rect -261 -704 -158 -696
rect -138 -704 61 -679
rect -261 -721 -185 -704
rect -166 -721 -158 -704
rect -261 -729 -158 -721
rect -261 -730 -163 -729
rect -138 -752 60 -723
rect -138 -783 -79 -752
rect -6 -783 60 -752
rect -261 -804 -164 -803
rect -261 -812 -158 -804
rect -138 -811 60 -783
rect -261 -829 -185 -812
rect -166 -829 -158 -812
rect -261 -837 -158 -829
rect -138 -860 60 -831
rect -138 -891 -76 -860
rect -4 -891 60 -860
rect -138 -920 60 -891
<< labels >>
rlabel locali 171 415 171 415 3 out
port 1 e
rlabel metal1 -122 518 -122 518 1 VDD
rlabel metal1 -261 443 -261 443 7 GND
rlabel metal1 -261 238 -261 238 7 A0
port 2 w
rlabel metal1 -260 133 -260 133 7 A1
port 3 w
rlabel metal1 -261 30 -261 30 7 A2
port 4 w
rlabel metal1 -261 -78 -261 -78 7 A3
port 5 w
rlabel metal1 -261 -188 -261 -188 7 A4
port 6 w
rlabel metal1 -261 -294 -261 -294 7 A5
port 7 w
rlabel metal1 -261 -401 -261 -401 7 A6
port 8 w
rlabel metal1 -261 -506 -261 -506 7 A7
port 9 w
rlabel metal1 -261 -608 -261 -608 7 A8
port 10 w
rlabel metal1 -261 -711 -261 -711 7 A9
port 11 w
rlabel metal1 -261 -821 -261 -821 7 A10
port 12 w
<< end >>
