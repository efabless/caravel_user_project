`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***
//***Module***
module parity_calculator #(
        parameter integer WORD_SIZE = 32,
        parameter integer ECCBITS = 7
    )
    (
        input  [WORD_SIZE - 1 : 0] data_to_register_i ,
        input  operate_i ,
        output [ECCBITS - 1 : 0] parity_bits_o ,
        output [WORD_SIZE - 1 : 0] data_to_register_o 
    );

//***Internal logic generated by compiler***  


//***Dumped Internal logic***
    assign  parity_bits_o[0] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[1] ^ data_to_register_i[3] ^ data_to_register_i[4]^ data_to_register_i[6]^ data_to_register_i[8]^ data_to_register_i[10]^ data_to_register_i[11]^ data_to_register_i[13]^ data_to_register_i[15]^ data_to_register_i[17]^ data_to_register_i[19]^ data_to_register_i[21]^ data_to_register_i[23] ^ data_to_register_i[25] ^ data_to_register_i[26]^ data_to_register_i[28]^ data_to_register_i[30] : 1'b0;
    assign  parity_bits_o[1] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[5]^ data_to_register_i[6]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[12]^ data_to_register_i[13]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[24] ^ data_to_register_i[25] ^ data_to_register_i[27]^ data_to_register_i[28]^ data_to_register_i[31] : 1'b0;
    assign  parity_bits_o[2] = operate_i ?  data_to_register_i[1] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24] ^ data_to_register_i[25] ^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31] : 1'b0;
    assign  parity_bits_o[3] = operate_i ?  data_to_register_i[4] ^ data_to_register_i[5] ^ data_to_register_i[6] ^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24] ^ data_to_register_i[25] : 1'b0;
    assign  parity_bits_o[4] = operate_i ?  data_to_register_i[11] ^ data_to_register_i[12] ^ data_to_register_i[13] ^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24]^ data_to_register_i[25]: 1'b0;
    assign  parity_bits_o[5] = operate_i ?  data_to_register_i[26] ^ data_to_register_i[27] ^ data_to_register_i[28] ^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31]: 1'b0;
    assign  parity_bits_o[6] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[1] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[4]^ data_to_register_i[5]^ data_to_register_i[6]^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[11]^ data_to_register_i[12]^ data_to_register_i[13]^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24]^ data_to_register_i[25]^ data_to_register_i[26]^ data_to_register_i[27]^ data_to_register_i[28]^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31]: 1'b0;
    assign  data_to_register_o = data_to_register_i;
    
//***Handcrafted Internal logic*** 
//TODO
endmodule
