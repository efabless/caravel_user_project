magic
tech sky130A
magscale 1 2
timestamp 1639940534
<< nwell >>
rect 786 330 1265 703
<< pwell >>
rect 1359 -264 2119 242
<< psubdiff >>
rect 1470 -94 1552 -68
rect 1470 -128 1492 -94
rect 1526 -128 1552 -94
rect 1470 -152 1552 -128
<< nsubdiff >>
rect 844 506 894 596
rect 828 504 900 506
rect 828 470 852 504
rect 886 470 900 504
rect 828 446 900 470
<< psubdiffcont >>
rect 1492 -128 1526 -94
<< nsubdiffcont >>
rect 852 470 886 504
<< locali >>
rect 844 648 930 682
rect 844 506 894 648
rect 828 504 900 506
rect 828 470 852 504
rect 886 470 900 504
rect 828 446 900 470
rect 842 330 954 342
rect 842 289 990 330
rect 842 206 900 289
rect 842 172 854 206
rect 888 172 900 206
rect 842 164 900 172
rect 1476 -68 1542 -16
rect 1470 -94 1552 -68
rect 1470 -128 1492 -94
rect 1526 -128 1552 -94
rect 1470 -152 1552 -128
rect 1600 -684 1602 -650
<< viali >>
rect 1864 528 1898 562
rect 1389 316 1423 350
rect 2978 260 3014 294
rect 854 172 888 206
rect 1931 -300 1965 -266
rect 2199 -310 2233 -276
rect 1723 -410 1757 -376
<< metal1 >>
rect 820 713 1609 714
rect 820 615 3077 713
rect 1852 562 1910 574
rect 820 528 1864 562
rect 1898 528 1910 562
rect 1852 516 1910 528
rect 1372 354 1440 362
rect 1372 350 1442 354
rect 1372 316 1389 350
rect 1423 340 1442 350
rect 1690 350 1766 354
rect 1690 340 1698 350
rect 1423 316 1698 340
rect 1372 308 1698 316
rect 1372 294 1438 308
rect 1686 298 1698 308
rect 1760 298 1766 350
rect 1686 294 1766 298
rect 2966 306 3080 308
rect 2966 254 2974 306
rect 3030 254 3080 306
rect 2966 248 3080 254
rect 840 208 900 216
rect 820 206 900 208
rect 820 172 854 206
rect 888 172 900 206
rect 820 160 900 172
rect 820 -51 3077 48
rect 2954 -92 3030 -84
rect 2954 -100 2968 -92
rect 2308 -136 2968 -100
rect 1920 -266 1974 -252
rect 2308 -258 2344 -136
rect 2954 -146 2968 -136
rect 3022 -146 3030 -92
rect 2954 -152 3030 -146
rect 1920 -270 1931 -266
rect 817 -300 1931 -270
rect 1965 -300 1974 -266
rect 817 -312 1974 -300
rect 2182 -276 2344 -258
rect 2182 -310 2199 -276
rect 2233 -310 2344 -276
rect 2182 -326 2344 -310
rect 1706 -362 1780 -356
rect 1706 -416 1712 -362
rect 1774 -416 1780 -362
rect 1706 -422 1780 -416
<< via1 >>
rect 1698 298 1760 350
rect 2974 294 3030 306
rect 2974 260 2978 294
rect 2978 260 3014 294
rect 3014 260 3030 294
rect 2974 254 3030 260
rect 2968 -146 3022 -92
rect 1712 -376 1774 -362
rect 1712 -410 1723 -376
rect 1723 -410 1757 -376
rect 1757 -410 1774 -376
rect 1712 -416 1774 -410
<< metal2 >>
rect 1692 350 1766 354
rect 1692 298 1698 350
rect 1760 298 1766 350
rect 1692 294 1766 298
rect 2966 306 3040 308
rect 1706 -356 1752 294
rect 2966 254 2974 306
rect 3030 254 3040 306
rect 2966 248 3040 254
rect 2966 -82 3022 248
rect 2958 -92 3030 -82
rect 2958 -146 2968 -92
rect 3022 -146 3030 -92
rect 2958 -156 3030 -146
rect 1706 -362 1780 -356
rect 1706 -416 1712 -362
rect 1774 -416 1780 -362
rect 1706 -422 1780 -416
use sky130_fd_sc_lp__dfrtp_1  sky130_fd_sc_lp__dfrtp_1_1 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 930 0 1 -1
box -38 -49 2150 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_1 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform -1 0 2274 0 -1 -1
box -38 -49 710 715
use sky130_fd_sc_lp__dfrtp_1  sky130_fd_sc_lp__dfrtp_1_0
timestamp 1626515395
transform 1 0 930 0 1 -1
box -38 -49 2150 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0
timestamp 1626515395
transform -1 0 2274 0 -1 -1
box -38 -49 710 715
use sky130_fd_sc_lp__dfrtp_1  sky130_fd_sc_lp__dfrtp_1_2
timestamp 1626515395
transform 1 0 930 0 1 -1
box -38 -49 2150 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_2
timestamp 1626515395
transform -1 0 2274 0 -1 -1
box -38 -49 710 715
use sky130_fd_sc_lp__dfrtp_1  sky130_fd_sc_lp__dfrtp_1_3
timestamp 1626515395
transform 1 0 930 0 1 -1
box -38 -49 2150 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_3
timestamp 1626515395
transform -1 0 2274 0 -1 -1
box -38 -49 710 715
<< end >>
