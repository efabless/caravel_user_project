magic
tech sky130A
timestamp 1640674630
<< locali >>
rect 3101 115 3142 126
rect 3101 98 3113 115
rect 3130 98 3142 115
rect 3101 82 3142 98
rect 3101 10 3142 21
rect 3101 -7 3113 10
rect 3130 -7 3142 10
rect 3101 -20 3142 -7
<< viali >>
rect 3113 98 3130 115
rect 3113 -7 3130 10
<< metal1 >>
rect -252 180 3179 201
rect -252 143 5 157
rect 186 143 3179 157
rect 3096 122 3148 127
rect 3096 107 3106 122
rect -252 93 4 107
rect 153 93 3106 107
rect 3138 107 3148 122
rect 3096 90 3106 93
rect 3138 93 3179 107
rect 3138 90 3148 93
rect 3096 76 3148 90
rect -252 46 7 60
rect 186 46 3179 60
rect -252 16 3179 21
rect -252 0 3107 16
rect 3101 -14 3107 0
rect 3136 0 3179 16
rect 3136 -14 3142 0
rect 3101 -20 3142 -14
<< via1 >>
rect 3106 115 3138 122
rect 3106 98 3113 115
rect 3113 98 3130 115
rect 3130 98 3138 115
rect 3106 90 3138 98
rect 3107 10 3136 16
rect 3107 -7 3113 10
rect 3113 -7 3130 10
rect 3130 -7 3136 10
rect 3107 -14 3136 -7
<< metal2 >>
rect 3096 122 3148 127
rect 3096 90 3106 122
rect 3138 90 3148 122
rect 3096 75 3148 90
rect 3101 16 3142 21
rect 3101 -14 3107 16
rect 3136 -14 3142 16
rect 3101 -20 3142 -14
<< via2 >>
rect 3106 90 3138 122
rect 3107 -14 3136 16
<< metal3 >>
rect 3096 122 3148 127
rect 3096 90 3106 122
rect 3138 90 3148 122
rect 3096 75 3148 90
rect 3096 16 3148 21
rect 3096 -14 3107 16
rect 3136 -14 3148 16
rect 3096 -30 3148 -14
<< via3 >>
rect 3106 90 3138 122
<< metal4 >>
rect 2967 515 3128 570
rect 3096 127 3128 515
rect 3096 122 3148 127
rect 3096 90 3106 122
rect 3138 90 3148 122
rect 3096 75 3148 90
use mimcap_8_32  mimcap_8_32_0
timestamp 1640667123
transform 1 0 8174 0 1 -475
box -8417 249 -5118 1077
use TG_min_dim  TG_min_dim_0
timestamp 1640671356
transform 1 0 78 0 1 33
box -78 -33 110 168
<< end >>
