* SPICE3 file created from asyn_rst_8_gray_counter.ext - technology: sky130A

.option scale=5000u

.subckt sky130_fd_sc_lp__xor2_1 A B VGND VNB VPB VPWR X a_293_367# a_42_367# a_297_69#
+ a_125_367#
X0 VPWR B a_293_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X1 a_297_69# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X2 a_125_367# B a_42_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X3 VGND a_42_367# X VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X4 a_42_367# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X5 X B a_297_69# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X6 a_293_367# a_42_367# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X7 a_293_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X8 VPWR A a_125_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X9 VGND A a_42_367# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
.ends

.subckt sky130_fd_sc_lp__and2_1 A B VGND VNB VPB VPWR X
X0 X a_92_131# VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X1 VGND B a_175_131# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X2 a_175_131# A a_92_131# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X3 a_92_131# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X4 X a_92_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X5 VPWR B a_92_131# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
.ends

.subckt sky130_fd_sc_lp__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q a_492_149# a_1467_419#
+ a_559_533# a_653_533# a_1417_133# a_196_462# a_1832_367# a_1593_133# a_1379_517#
+ a_695_375# a_304_533# a_27_114# a_803_149# a_1247_89# a_875_149#
X0 a_492_149# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X1 VGND a_1467_419# a_1417_133# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X2 a_803_149# a_196_462# a_559_533# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X3 a_1379_517# a_196_462# a_1247_89# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X4 VPWR a_695_375# a_653_533# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X5 a_559_533# a_27_114# a_304_533# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X6 a_1417_133# a_27_114# a_1247_89# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X7 a_1467_419# a_1247_89# a_1593_133# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X8 a_695_375# a_559_533# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=168 l=30
X9 a_559_533# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X10 a_1593_133# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X11 VPWR RESET_B a_304_533# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X12 a_695_375# a_559_533# VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=128 l=30
X13 a_653_533# a_27_114# a_559_533# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X14 a_196_462# a_27_114# VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X15 a_1247_89# a_27_114# a_695_375# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=168 l=30
X16 VGND RESET_B a_875_149# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X17 a_196_462# a_27_114# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=128 l=30
X18 a_304_533# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X19 VPWR CLK a_27_114# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=128 l=30
X20 VPWR a_1247_89# a_1467_419# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X21 Q a_1832_367# VGND VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=168 l=30
X22 a_1467_419# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X23 a_304_533# D a_492_149# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X24 a_875_149# a_695_375# a_803_149# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X25 VGND a_1247_89# a_1832_367# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X26 a_559_533# a_196_462# a_304_533# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X27 VPWR a_1467_419# a_1379_517# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=84 l=30
X28 VPWR a_1247_89# a_1832_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=128 l=30
X29 VGND CLK a_27_114# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=84 l=30
X30 Q a_1832_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=252 l=30
X31 a_1247_89# a_196_462# a_695_375# VNB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=128 l=30
.ends

.subckt T_flip_flop sky130_fd_sc_lp__xor2_1_3/A sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VPB sky130_fd_sc_lp__dfrtp_1_3/RESET_B
+ sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__dfrtp_1_3/CLK
Xsky130_fd_sc_lp__dfrtp_1_3 sky130_fd_sc_lp__dfrtp_1_3/CLK sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB
+ sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__dfrtp_1_3/a_492_149# sky130_fd_sc_lp__dfrtp_1_3/a_1467_419# sky130_fd_sc_lp__dfrtp_1_3/a_559_533#
+ sky130_fd_sc_lp__dfrtp_1_3/a_653_533# sky130_fd_sc_lp__dfrtp_1_3/a_1417_133# sky130_fd_sc_lp__dfrtp_1_3/a_196_462#
+ sky130_fd_sc_lp__dfrtp_1_3/a_1832_367# sky130_fd_sc_lp__dfrtp_1_3/a_1593_133# sky130_fd_sc_lp__dfrtp_1_3/a_1379_517#
+ sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__dfrtp_1_3/a_304_533# sky130_fd_sc_lp__dfrtp_1_3/a_27_114#
+ sky130_fd_sc_lp__dfrtp_1_3/a_803_149# sky130_fd_sc_lp__dfrtp_1_3/a_1247_89# sky130_fd_sc_lp__dfrtp_1_3/a_875_149#
+ sky130_fd_sc_lp__dfrtp_1
Xsky130_fd_sc_lp__xor2_1_0 sky130_fd_sc_lp__xor2_1_3/A sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VPB
+ sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__xor2_1_3/X sky130_fd_sc_lp__xor2_1_3/a_293_367#
+ sky130_fd_sc_lp__xor2_1_3/a_42_367# sky130_fd_sc_lp__xor2_1_3/a_297_69# sky130_fd_sc_lp__xor2_1_3/a_125_367#
+ sky130_fd_sc_lp__xor2_1
Xsky130_fd_sc_lp__xor2_1_1 sky130_fd_sc_lp__xor2_1_3/A sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VPB
+ sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__xor2_1_3/X sky130_fd_sc_lp__xor2_1_3/a_293_367#
+ sky130_fd_sc_lp__xor2_1_3/a_42_367# sky130_fd_sc_lp__xor2_1_3/a_297_69# sky130_fd_sc_lp__xor2_1_3/a_125_367#
+ sky130_fd_sc_lp__xor2_1
Xsky130_fd_sc_lp__xor2_1_2 sky130_fd_sc_lp__xor2_1_3/A sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VPB
+ sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__xor2_1_3/X sky130_fd_sc_lp__xor2_1_3/a_293_367#
+ sky130_fd_sc_lp__xor2_1_3/a_42_367# sky130_fd_sc_lp__xor2_1_3/a_297_69# sky130_fd_sc_lp__xor2_1_3/a_125_367#
+ sky130_fd_sc_lp__xor2_1
Xsky130_fd_sc_lp__xor2_1_3 sky130_fd_sc_lp__xor2_1_3/A sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VPB
+ sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__xor2_1_3/X sky130_fd_sc_lp__xor2_1_3/a_293_367#
+ sky130_fd_sc_lp__xor2_1_3/a_42_367# sky130_fd_sc_lp__xor2_1_3/a_297_69# sky130_fd_sc_lp__xor2_1_3/a_125_367#
+ sky130_fd_sc_lp__xor2_1
Xsky130_fd_sc_lp__dfrtp_1_0 sky130_fd_sc_lp__dfrtp_1_3/CLK sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB
+ sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__dfrtp_1_3/a_492_149# sky130_fd_sc_lp__dfrtp_1_3/a_1467_419# sky130_fd_sc_lp__dfrtp_1_3/a_559_533#
+ sky130_fd_sc_lp__dfrtp_1_3/a_653_533# sky130_fd_sc_lp__dfrtp_1_3/a_1417_133# sky130_fd_sc_lp__dfrtp_1_3/a_196_462#
+ sky130_fd_sc_lp__dfrtp_1_3/a_1832_367# sky130_fd_sc_lp__dfrtp_1_3/a_1593_133# sky130_fd_sc_lp__dfrtp_1_3/a_1379_517#
+ sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__dfrtp_1_3/a_304_533# sky130_fd_sc_lp__dfrtp_1_3/a_27_114#
+ sky130_fd_sc_lp__dfrtp_1_3/a_803_149# sky130_fd_sc_lp__dfrtp_1_3/a_1247_89# sky130_fd_sc_lp__dfrtp_1_3/a_875_149#
+ sky130_fd_sc_lp__dfrtp_1
Xsky130_fd_sc_lp__dfrtp_1_1 sky130_fd_sc_lp__dfrtp_1_3/CLK sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB
+ sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__dfrtp_1_3/a_492_149# sky130_fd_sc_lp__dfrtp_1_3/a_1467_419# sky130_fd_sc_lp__dfrtp_1_3/a_559_533#
+ sky130_fd_sc_lp__dfrtp_1_3/a_653_533# sky130_fd_sc_lp__dfrtp_1_3/a_1417_133# sky130_fd_sc_lp__dfrtp_1_3/a_196_462#
+ sky130_fd_sc_lp__dfrtp_1_3/a_1832_367# sky130_fd_sc_lp__dfrtp_1_3/a_1593_133# sky130_fd_sc_lp__dfrtp_1_3/a_1379_517#
+ sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__dfrtp_1_3/a_304_533# sky130_fd_sc_lp__dfrtp_1_3/a_27_114#
+ sky130_fd_sc_lp__dfrtp_1_3/a_803_149# sky130_fd_sc_lp__dfrtp_1_3/a_1247_89# sky130_fd_sc_lp__dfrtp_1_3/a_875_149#
+ sky130_fd_sc_lp__dfrtp_1
Xsky130_fd_sc_lp__dfrtp_1_2 sky130_fd_sc_lp__dfrtp_1_3/CLK sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_3/VNB sky130_fd_sc_lp__xor2_1_3/VNB
+ sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/B
+ sky130_fd_sc_lp__dfrtp_1_3/a_492_149# sky130_fd_sc_lp__dfrtp_1_3/a_1467_419# sky130_fd_sc_lp__dfrtp_1_3/a_559_533#
+ sky130_fd_sc_lp__dfrtp_1_3/a_653_533# sky130_fd_sc_lp__dfrtp_1_3/a_1417_133# sky130_fd_sc_lp__dfrtp_1_3/a_196_462#
+ sky130_fd_sc_lp__dfrtp_1_3/a_1832_367# sky130_fd_sc_lp__dfrtp_1_3/a_1593_133# sky130_fd_sc_lp__dfrtp_1_3/a_1379_517#
+ sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__dfrtp_1_3/a_304_533# sky130_fd_sc_lp__dfrtp_1_3/a_27_114#
+ sky130_fd_sc_lp__dfrtp_1_3/a_803_149# sky130_fd_sc_lp__dfrtp_1_3/a_1247_89# sky130_fd_sc_lp__dfrtp_1_3/a_875_149#
+ sky130_fd_sc_lp__dfrtp_1
C0 sky130_fd_sc_lp__dfrtp_1_3/a_1247_89# sky130_fd_sc_lp__xor2_1_3/VNB -2.03fF
C1 sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__xor2_1_3/VNB 2.41fF
C2 sky130_fd_sc_lp__dfrtp_1_3/a_196_462# sky130_fd_sc_lp__xor2_1_3/VNB 3.49fF
C3 sky130_fd_sc_lp__xor2_1_3/VPWR sky130_fd_sc_lp__xor2_1_3/VNB 2.17fF
C4 sky130_fd_sc_lp__xor2_1_3/B sky130_fd_sc_lp__xor2_1_3/VNB 3.19fF
C5 sky130_fd_sc_lp__xor2_1_3/VPB sky130_fd_sc_lp__xor2_1_3/VNB 2.70fF
C6 sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_3/VNB -3.79fF
C7 sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_3/VNB 10.00fF
.ends

.subckt asyn_rst_counter_cell T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/VPB T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/RESET_B
+ sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__and2_1_0/B sky130_fd_sc_lp__xor2_1_0/VPB
+ sky130_fd_sc_lp__xor2_1_0/VPWR sky130_fd_sc_lp__xor2_1_0/A sky130_fd_sc_lp__xor2_1_0/B
+ T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/CLK sky130_fd_sc_lp__and2_1_0/X
Xsky130_fd_sc_lp__xor2_1_0 sky130_fd_sc_lp__xor2_1_0/A sky130_fd_sc_lp__xor2_1_0/B
+ sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__xor2_1_0/VPB
+ sky130_fd_sc_lp__xor2_1_0/VPWR sky130_fd_sc_lp__xor2_1_0/X sky130_fd_sc_lp__xor2_1_0/a_293_367#
+ sky130_fd_sc_lp__xor2_1_0/a_42_367# sky130_fd_sc_lp__xor2_1_0/a_297_69# sky130_fd_sc_lp__xor2_1_0/a_125_367#
+ sky130_fd_sc_lp__xor2_1
Xsky130_fd_sc_lp__and2_1_0 sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__xor2_1_0/VPB
+ sky130_fd_sc_lp__xor2_1_0/VPWR sky130_fd_sc_lp__and2_1_0/X sky130_fd_sc_lp__and2_1
XT_flip_flop_0 sky130_fd_sc_lp__and2_1_0/B T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/VPB
+ sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__xor2_1_0/VNB sky130_fd_sc_lp__xor2_1_0/VPB
+ T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_0/VPWR
+ T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/CLK T_flip_flop
C0 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# sky130_fd_sc_lp__xor2_1_0/VNB 2.21fF
C1 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# sky130_fd_sc_lp__xor2_1_0/VNB 2.57fF
C2 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# sky130_fd_sc_lp__xor2_1_0/VNB 5.90fF
C3 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# sky130_fd_sc_lp__xor2_1_0/VNB 4.23fF
C4 sky130_fd_sc_lp__xor2_1_0/VPWR sky130_fd_sc_lp__xor2_1_0/VNB 3.77fF
C5 sky130_fd_sc_lp__and2_1_0/B sky130_fd_sc_lp__xor2_1_0/VNB 2.14fF
C6 sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__xor2_1_0/VNB 6.05fF
C7 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/RESET_B sky130_fd_sc_lp__xor2_1_0/VNB -2.74fF
C8 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/VPB sky130_fd_sc_lp__xor2_1_0/VNB 10.24fF
C9 sky130_fd_sc_lp__xor2_1_0/VPB sky130_fd_sc_lp__xor2_1_0/VNB 5.61fF
.ends

.subckt asyn_rst_8_gray_counter RSTB CLK Vdd gnd
Xasyn_rst_counter_cell_1 Vdd RSTB gnd asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
Xasyn_rst_counter_cell_2 Vdd RSTB gnd asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
Xasyn_rst_counter_cell_3 Vdd RSTB gnd asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
Xasyn_rst_counter_cell_4 Vdd RSTB gnd asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
Xasyn_rst_counter_cell_5 Vdd RSTB gnd asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
Xasyn_rst_counter_cell_6 Vdd RSTB gnd asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B
+ CLK T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A asyn_rst_counter_cell
XT_flip_flop_0 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B
+ gnd Vdd RSTB Vdd CLK T_flip_flop
Xasyn_rst_counter_cell_0 Vdd RSTB gnd asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B
+ Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B
+ CLK asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B asyn_rst_counter_cell
C0 RSTB CLK 11.27fF
C1 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C2 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C3 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C4 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C5 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B gnd 2.02fF
C6 asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd 4.57fF
C7 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.02fF
C8 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C9 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C10 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C11 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A gnd 2.28fF
C12 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd 4.10fF
C13 Vdd gnd 176.79fF
C14 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.02fF
C15 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C16 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C17 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C18 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C19 asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
C20 CLK gnd 17.32fF
C21 RSTB gnd -17.29fF
C22 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C23 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C24 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C25 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C26 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C27 asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
C28 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C29 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C30 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C31 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C32 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C33 asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
C34 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C35 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C36 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C37 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C38 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C39 asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
C40 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C41 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C42 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C43 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C44 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C45 asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
C46 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.12fF
C47 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.57fF
C48 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 5.90fF
C49 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.23fF
C50 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B gnd 2.45fF
C51 asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd 5.40fF
.ends

