VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_4kbyte_1rw_64x512_8
   CLASS BLOCK ;
   SIZE 828.62 BY 339.02 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 0.0 178.54 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  184.28 0.0 184.66 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.72 0.0 190.1 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.52 0.0 196.9 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.64 0.0 203.02 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 0.0 207.78 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.2 0.0 214.58 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  219.64 0.0 220.02 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.08 0.0 225.46 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  236.64 0.0 237.02 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.44 0.0 243.82 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.32 0.0 254.7 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 0.0 260.14 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.56 0.0 283.94 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 0.0 289.38 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.8 0.0 296.18 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  301.24 0.0 301.62 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.68 0.0 307.06 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 0.0 313.18 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  318.24 0.0 318.62 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  325.04 0.0 325.42 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  331.16 0.0 331.54 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  335.92 0.0 336.3 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  342.04 0.0 342.42 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  347.48 0.0 347.86 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  354.28 0.0 354.66 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  359.72 0.0 360.1 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  365.16 0.0 365.54 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 0.0 372.34 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  377.4 0.0 377.78 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  382.84 0.0 383.22 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  388.28 0.0 388.66 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  394.4 0.0 394.78 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  401.2 0.0 401.58 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  412.08 0.0 412.46 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  417.52 0.0 417.9 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  423.64 0.0 424.02 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  430.44 0.0 430.82 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  435.88 0.0 436.26 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  441.32 0.0 441.7 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  446.76 0.0 447.14 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  453.56 0.0 453.94 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  459.0 0.0 459.38 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  464.44 0.0 464.82 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  471.24 0.0 471.62 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  476.0 0.0 476.38 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  482.8 0.0 483.18 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  488.24 0.0 488.62 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  493.68 0.0 494.06 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  499.12 0.0 499.5 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  505.24 0.0 505.62 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  512.04 0.0 512.42 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  517.48 0.0 517.86 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  522.92 0.0 523.3 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  529.72 0.0 530.1 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  535.16 0.0 535.54 1.06 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  540.6 0.0 540.98 1.06 ;
      END
   END din0[64]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.12 0.0 108.5 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  114.92 0.0 115.3 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.08 1.06 157.46 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 166.6 1.06 166.98 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 172.04 1.06 172.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 180.2 1.06 180.58 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 185.64 1.06 186.02 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 194.48 1.06 194.86 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 200.6 1.06 200.98 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 208.76 1.06 209.14 ;
      END
   END addr0[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 54.4 1.06 54.78 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 63.24 1.06 63.62 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 55.08 1.06 55.46 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  120.36 0.0 120.74 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.8 0.0 126.18 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.6 0.0 132.98 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.04 0.0 138.42 1.06 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 1.06 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.92 0.0 149.3 1.06 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  155.04 0.0 155.42 1.06 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 0.0 160.86 1.06 ;
      END
   END wmask0[7]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  546.04 0.0 546.42 1.06 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 0.0 182.62 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 0.0 211.86 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 0.0 243.14 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  281.52 0.0 281.9 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.76 0.0 311.14 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.32 0.0 322.7 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 0.0 330.86 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 0.0 343.1 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  351.56 0.0 351.94 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  362.44 0.0 362.82 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  372.64 0.0 373.02 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  380.8 0.0 381.18 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  392.36 0.0 392.74 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  402.56 0.0 402.94 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  410.04 0.0 410.42 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  421.6 0.0 421.98 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  432.48 0.0 432.86 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  442.68 0.0 443.06 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  452.88 0.0 453.26 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  462.4 0.0 462.78 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  472.6 0.0 472.98 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  482.12 0.0 482.5 1.06 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  490.96 0.0 491.34 1.06 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  502.52 0.0 502.9 1.06 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  512.72 0.0 513.1 1.06 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  520.88 0.0 521.26 1.06 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  532.44 0.0 532.82 1.06 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  542.64 0.0 543.02 1.06 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  552.84 0.0 553.22 1.06 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  562.36 0.0 562.74 1.06 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  571.2 0.0 571.58 1.06 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  582.08 0.0 582.46 1.06 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  592.28 0.0 592.66 1.06 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  602.48 0.0 602.86 1.06 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  612.68 0.0 613.06 1.06 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  622.88 0.0 623.26 1.06 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  632.4 0.0 632.78 1.06 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  642.6 0.0 642.98 1.06 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  651.44 0.0 651.82 1.06 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  662.32 0.0 662.7 1.06 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  672.52 0.0 672.9 1.06 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  682.72 0.0 683.1 1.06 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  692.24 0.0 692.62 1.06 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  702.44 0.0 702.82 1.06 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  712.64 0.0 713.02 1.06 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  722.16 0.0 722.54 1.06 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  731.0 0.0 731.38 1.06 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  742.56 0.0 742.94 1.06 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  752.76 0.0 753.14 1.06 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 83.64 828.62 84.02 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 78.88 828.62 79.26 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 82.96 828.62 83.34 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 76.84 828.62 77.22 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 82.28 828.62 82.66 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  827.56 80.24 828.62 80.62 ;
      END
   END dout0[64]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  822.12 4.76 823.86 335.62 ;
         LAYER met3 ;
         RECT  4.76 4.76 823.86 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 335.62 ;
         LAYER met3 ;
         RECT  4.76 333.88 823.86 335.62 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  1.36 337.28 827.26 339.02 ;
         LAYER met4 ;
         RECT  825.52 1.36 827.26 339.02 ;
         LAYER met3 ;
         RECT  1.36 1.36 827.26 3.1 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 339.02 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 828.0 338.4 ;
   LAYER  met2 ;
      RECT  0.62 0.62 828.0 338.4 ;
   LAYER  met3 ;
      RECT  1.66 156.48 828.0 158.06 ;
      RECT  0.62 158.06 1.66 166.0 ;
      RECT  0.62 167.58 1.66 171.44 ;
      RECT  0.62 173.02 1.66 179.6 ;
      RECT  0.62 181.18 1.66 185.04 ;
      RECT  0.62 186.62 1.66 193.88 ;
      RECT  0.62 195.46 1.66 200.0 ;
      RECT  0.62 201.58 1.66 208.16 ;
      RECT  0.62 64.22 1.66 156.48 ;
      RECT  0.62 56.06 1.66 62.64 ;
      RECT  1.66 83.04 826.96 84.62 ;
      RECT  1.66 84.62 826.96 156.48 ;
      RECT  826.96 84.62 828.0 156.48 ;
      RECT  826.96 77.82 828.0 78.28 ;
      RECT  826.96 81.22 828.0 81.68 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 83.04 ;
      RECT  4.16 7.1 824.46 83.04 ;
      RECT  824.46 4.16 826.96 7.1 ;
      RECT  824.46 7.1 826.96 83.04 ;
      RECT  1.66 158.06 4.16 333.28 ;
      RECT  1.66 333.28 4.16 336.22 ;
      RECT  4.16 158.06 824.46 333.28 ;
      RECT  824.46 158.06 828.0 333.28 ;
      RECT  824.46 333.28 828.0 336.22 ;
      RECT  0.62 209.74 0.76 336.68 ;
      RECT  0.62 336.68 0.76 338.4 ;
      RECT  0.76 209.74 1.66 336.68 ;
      RECT  1.66 336.22 4.16 336.68 ;
      RECT  4.16 336.22 824.46 336.68 ;
      RECT  824.46 336.22 827.86 336.68 ;
      RECT  827.86 336.22 828.0 336.68 ;
      RECT  827.86 336.68 828.0 338.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 53.8 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 53.8 ;
      RECT  826.96 0.62 827.86 0.76 ;
      RECT  826.96 3.7 827.86 76.24 ;
      RECT  827.86 0.62 828.0 0.76 ;
      RECT  827.86 0.76 828.0 3.7 ;
      RECT  827.86 3.7 828.0 76.24 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 824.46 0.76 ;
      RECT  4.16 3.7 824.46 4.16 ;
      RECT  824.46 0.62 826.96 0.76 ;
      RECT  824.46 3.7 826.96 4.16 ;
   LAYER  met4 ;
      RECT  166.68 1.66 168.26 338.4 ;
      RECT  173.7 0.62 177.56 1.66 ;
      RECT  185.26 0.62 189.12 1.66 ;
      RECT  203.62 0.62 206.8 1.66 ;
      RECT  215.18 0.62 219.04 1.66 ;
      RECT  226.06 0.62 231.28 1.66 ;
      RECT  244.42 0.62 248.28 1.66 ;
      RECT  255.3 0.62 259.16 1.66 ;
      RECT  273.66 0.62 277.52 1.66 ;
      RECT  284.54 0.62 288.4 1.66 ;
      RECT  296.78 0.62 300.64 1.66 ;
      RECT  313.78 0.62 317.64 1.66 ;
      RECT  332.14 0.62 335.32 1.66 ;
      RECT  336.9 0.62 341.44 1.66 ;
      RECT  355.26 0.62 359.12 1.66 ;
      RECT  366.14 0.62 371.36 1.66 ;
      RECT  383.82 0.62 387.68 1.66 ;
      RECT  395.38 0.62 400.6 1.66 ;
      RECT  413.06 0.62 416.92 1.66 ;
      RECT  424.62 0.62 429.84 1.66 ;
      RECT  436.86 0.62 440.72 1.66 ;
      RECT  454.54 0.62 458.4 1.66 ;
      RECT  465.42 0.62 470.64 1.66 ;
      RECT  483.78 0.62 487.64 1.66 ;
      RECT  494.66 0.62 498.52 1.66 ;
      RECT  506.22 0.62 511.44 1.66 ;
      RECT  523.9 0.62 529.12 1.66 ;
      RECT  536.14 0.62 540.0 1.66 ;
      RECT  109.1 0.62 114.32 1.66 ;
      RECT  115.9 0.62 119.76 1.66 ;
      RECT  121.34 0.62 125.2 1.66 ;
      RECT  126.78 0.62 132.0 1.66 ;
      RECT  133.58 0.62 137.44 1.66 ;
      RECT  139.02 0.62 142.88 1.66 ;
      RECT  144.46 0.62 148.32 1.66 ;
      RECT  149.9 0.62 154.44 1.66 ;
      RECT  156.02 0.62 159.88 1.66 ;
      RECT  161.46 0.62 166.68 1.66 ;
      RECT  168.26 0.62 170.08 1.66 ;
      RECT  171.66 0.62 172.12 1.66 ;
      RECT  179.14 0.62 181.64 1.66 ;
      RECT  183.22 0.62 183.68 1.66 ;
      RECT  190.7 0.62 191.84 1.66 ;
      RECT  193.42 0.62 195.92 1.66 ;
      RECT  197.5 0.62 201.36 1.66 ;
      RECT  208.38 0.62 210.88 1.66 ;
      RECT  212.46 0.62 213.6 1.66 ;
      RECT  220.62 0.62 221.76 1.66 ;
      RECT  223.34 0.62 224.48 1.66 ;
      RECT  233.54 0.62 236.04 1.66 ;
      RECT  237.62 0.62 242.16 1.66 ;
      RECT  249.86 0.62 250.32 1.66 ;
      RECT  251.9 0.62 253.72 1.66 ;
      RECT  260.74 0.62 261.88 1.66 ;
      RECT  263.46 0.62 265.28 1.66 ;
      RECT  266.86 0.62 271.4 1.66 ;
      RECT  279.1 0.62 280.92 1.66 ;
      RECT  282.5 0.62 282.96 1.66 ;
      RECT  289.98 0.62 291.8 1.66 ;
      RECT  293.38 0.62 295.2 1.66 ;
      RECT  303.58 0.62 306.08 1.66 ;
      RECT  307.66 0.62 310.16 1.66 ;
      RECT  311.74 0.62 312.2 1.66 ;
      RECT  319.22 0.62 321.72 1.66 ;
      RECT  323.3 0.62 324.44 1.66 ;
      RECT  326.02 0.62 329.88 1.66 ;
      RECT  343.7 0.62 346.88 1.66 ;
      RECT  348.46 0.62 350.96 1.66 ;
      RECT  352.54 0.62 353.68 1.66 ;
      RECT  360.7 0.62 361.84 1.66 ;
      RECT  363.42 0.62 364.56 1.66 ;
      RECT  373.62 0.62 376.8 1.66 ;
      RECT  378.38 0.62 380.2 1.66 ;
      RECT  381.78 0.62 382.24 1.66 ;
      RECT  389.26 0.62 391.76 1.66 ;
      RECT  393.34 0.62 393.8 1.66 ;
      RECT  403.54 0.62 406.04 1.66 ;
      RECT  407.62 0.62 409.44 1.66 ;
      RECT  411.02 0.62 411.48 1.66 ;
      RECT  418.5 0.62 421.0 1.66 ;
      RECT  422.58 0.62 423.04 1.66 ;
      RECT  431.42 0.62 431.88 1.66 ;
      RECT  433.46 0.62 435.28 1.66 ;
      RECT  443.66 0.62 446.16 1.66 ;
      RECT  447.74 0.62 452.28 1.66 ;
      RECT  459.98 0.62 461.8 1.66 ;
      RECT  463.38 0.62 463.84 1.66 ;
      RECT  473.58 0.62 475.4 1.66 ;
      RECT  476.98 0.62 481.52 1.66 ;
      RECT  489.22 0.62 490.36 1.66 ;
      RECT  491.94 0.62 493.08 1.66 ;
      RECT  500.1 0.62 501.92 1.66 ;
      RECT  503.5 0.62 504.64 1.66 ;
      RECT  513.7 0.62 516.88 1.66 ;
      RECT  518.46 0.62 520.28 1.66 ;
      RECT  521.86 0.62 522.32 1.66 ;
      RECT  530.7 0.62 531.84 1.66 ;
      RECT  533.42 0.62 534.56 1.66 ;
      RECT  541.58 0.62 542.04 1.66 ;
      RECT  543.62 0.62 545.44 1.66 ;
      RECT  547.02 0.62 552.24 1.66 ;
      RECT  553.82 0.62 561.76 1.66 ;
      RECT  563.34 0.62 570.6 1.66 ;
      RECT  572.18 0.62 581.48 1.66 ;
      RECT  583.06 0.62 591.68 1.66 ;
      RECT  593.26 0.62 601.88 1.66 ;
      RECT  603.46 0.62 612.08 1.66 ;
      RECT  613.66 0.62 622.28 1.66 ;
      RECT  623.86 0.62 631.8 1.66 ;
      RECT  633.38 0.62 642.0 1.66 ;
      RECT  643.58 0.62 650.84 1.66 ;
      RECT  652.42 0.62 661.72 1.66 ;
      RECT  663.3 0.62 671.92 1.66 ;
      RECT  673.5 0.62 682.12 1.66 ;
      RECT  683.7 0.62 691.64 1.66 ;
      RECT  693.22 0.62 701.84 1.66 ;
      RECT  703.42 0.62 712.04 1.66 ;
      RECT  713.62 0.62 721.56 1.66 ;
      RECT  723.14 0.62 730.4 1.66 ;
      RECT  731.98 0.62 741.96 1.66 ;
      RECT  743.54 0.62 752.16 1.66 ;
      RECT  168.26 1.66 821.52 4.16 ;
      RECT  168.26 4.16 821.52 336.22 ;
      RECT  168.26 336.22 821.52 338.4 ;
      RECT  821.52 1.66 824.46 4.16 ;
      RECT  821.52 336.22 824.46 338.4 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 336.22 7.1 338.4 ;
      RECT  7.1 1.66 166.68 4.16 ;
      RECT  7.1 4.16 166.68 336.22 ;
      RECT  7.1 336.22 166.68 338.4 ;
      RECT  753.74 0.62 824.92 0.76 ;
      RECT  753.74 0.76 824.92 1.66 ;
      RECT  824.92 0.62 827.86 0.76 ;
      RECT  827.86 0.62 828.0 0.76 ;
      RECT  827.86 0.76 828.0 1.66 ;
      RECT  824.46 1.66 824.92 4.16 ;
      RECT  827.86 1.66 828.0 4.16 ;
      RECT  824.46 4.16 824.92 336.22 ;
      RECT  827.86 4.16 828.0 336.22 ;
      RECT  824.46 336.22 824.92 338.4 ;
      RECT  827.86 336.22 828.0 338.4 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 107.52 0.76 ;
      RECT  3.7 0.76 107.52 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 336.22 ;
      RECT  3.7 4.16 4.16 336.22 ;
      RECT  0.62 336.22 0.76 338.4 ;
      RECT  3.7 336.22 4.16 338.4 ;
   END
END    sky130_sram_4kbyte_1rw_64x512_8
END    LIBRARY
