magic
tech sky130A
magscale 1 2
timestamp 1641166894
<< nwell >>
rect 142 10576 3292 10760
rect 2066 10374 2924 10576
rect 5365 10548 7124 10760
rect 5365 10530 5448 10548
rect 6748 10532 7124 10548
rect 5410 10482 5448 10530
rect 6750 10482 7124 10532
rect 2888 9712 2908 9912
rect 1769 9042 3005 9712
rect 1769 7710 2917 8380
rect 1769 6378 2939 7048
rect 1769 5046 2993 5716
rect 1769 3714 2929 4384
rect 1769 2382 3005 3052
rect 1769 1118 2965 1720
rect 5287 1272 7102 1354
rect 3035 1118 4654 1272
rect 4806 1118 7102 1272
rect 1769 1052 7102 1118
rect 1769 1050 4654 1052
rect 3035 694 4654 1050
<< locali >>
rect 2449 10738 5284 10739
rect 2448 10681 5284 10738
rect 2448 9898 2504 10681
rect 2538 10580 4444 10640
rect 2448 9674 2500 9898
rect 2448 9640 2456 9674
rect 2490 9640 2500 9674
rect 2448 9630 2500 9640
rect 2538 7008 2598 10580
rect 3524 10434 3542 10442
rect 2538 6974 2552 7008
rect 2586 6974 2598 7008
rect 2538 6966 2598 6974
rect 2640 10370 3542 10434
rect 4384 10370 4444 10580
rect 5226 10370 5284 10681
rect 7551 10522 7737 10588
rect 2640 4344 2704 10370
rect 5940 10228 5992 10242
rect 5940 10190 5952 10228
rect 5986 10190 5992 10228
rect 5940 10172 5992 10190
rect 5944 9634 5992 10172
rect 6356 10006 6414 10024
rect 6356 9972 6366 10006
rect 6404 9972 6414 10006
rect 6356 9956 6414 9972
rect 5944 9620 5984 9634
rect 6020 9516 6104 9524
rect 6226 9516 6306 9524
rect 6020 9510 6306 9516
rect 6020 9472 6256 9510
rect 6290 9472 6306 9510
rect 6020 9466 6306 9472
rect 6020 9460 6104 9466
rect 6226 9460 6306 9466
rect 5952 9268 5992 9340
rect 6356 9268 6396 9956
rect 6432 9800 6488 9818
rect 6432 9766 6440 9800
rect 6478 9766 6488 9800
rect 6432 9748 6488 9766
rect 5952 9228 6396 9268
rect 6434 8956 6474 9748
rect 6514 9584 6568 9604
rect 6514 9550 6522 9584
rect 6560 9550 6568 9584
rect 6514 9534 6568 9550
rect 5950 8916 6474 8956
rect 5950 8842 5990 8916
rect 6018 8716 6102 8726
rect 6224 8716 6306 8726
rect 6018 8706 6306 8716
rect 6018 8672 6254 8706
rect 6288 8672 6306 8706
rect 6018 8666 6306 8672
rect 6018 8656 6102 8666
rect 6224 8656 6306 8666
rect 5950 8448 5990 8540
rect 6516 8448 6556 9534
rect 5950 8408 6556 8448
rect 6598 9364 6650 9384
rect 6598 9330 6606 9364
rect 6644 9330 6650 9364
rect 6598 9314 6650 9330
rect 2640 4310 2654 4344
rect 2688 4310 2704 4344
rect 2640 4302 2704 4310
rect 2744 8340 2800 8350
rect 2744 8306 2756 8340
rect 2790 8306 2800 8340
rect 2660 1680 2708 1690
rect 2660 1646 2664 1680
rect 2698 1646 2708 1680
rect 2660 1072 2708 1646
rect 2744 1166 2800 8306
rect 6598 8158 6638 9314
rect 6672 9152 6720 9172
rect 6672 9118 6678 9152
rect 6716 9118 6720 9152
rect 6672 9104 6720 9118
rect 5950 8118 6638 8158
rect 5950 8042 5990 8118
rect 6018 7910 6102 7922
rect 6224 7910 6306 7922
rect 6018 7908 6306 7910
rect 6018 7874 6254 7908
rect 6288 7874 6306 7908
rect 6018 7868 6306 7874
rect 6018 7858 6102 7868
rect 6224 7858 6306 7868
rect 5950 7658 5990 7740
rect 6674 7658 6714 9104
rect 5950 7618 6714 7658
rect 6448 7358 6516 7368
rect 6448 7352 6464 7358
rect 5948 7320 6464 7352
rect 6498 7320 6516 7358
rect 5948 7312 6516 7320
rect 5948 7236 5988 7312
rect 6016 7116 6100 7122
rect 6222 7116 6306 7122
rect 6016 7108 6306 7116
rect 6016 7074 6254 7108
rect 6288 7074 6306 7108
rect 6016 7066 6306 7074
rect 6016 7058 6100 7066
rect 6222 7058 6306 7066
rect 5948 6864 5988 6942
rect 6570 6870 6638 6888
rect 6570 6864 6586 6870
rect 5948 6836 6586 6864
rect 6620 6836 6638 6870
rect 5948 6824 6638 6836
rect 6668 6540 6736 6554
rect 6668 6534 6686 6540
rect 5950 6506 6686 6534
rect 6720 6506 6736 6540
rect 5950 6494 6736 6506
rect 5950 6432 5990 6494
rect 6018 6316 6102 6330
rect 6224 6316 6306 6330
rect 6018 6310 6306 6316
rect 6018 6276 6256 6310
rect 6290 6276 6306 6310
rect 6018 6266 6306 6276
rect 6018 6258 6102 6266
rect 6224 6258 6306 6266
rect 5950 6086 5990 6140
rect 5950 6084 6626 6086
rect 5950 6070 6630 6084
rect 5950 6046 6576 6070
rect 6558 6036 6576 6046
rect 6610 6036 6630 6070
rect 6558 6024 6630 6036
rect 6768 5764 6836 5780
rect 6768 5756 6786 5764
rect 5946 5730 6786 5756
rect 6820 5730 6836 5764
rect 5946 5716 6836 5730
rect 2834 5678 2882 5686
rect 2834 5644 2842 5678
rect 2876 5644 2882 5678
rect 2834 1260 2882 5644
rect 5946 5642 5986 5716
rect 6014 5516 6098 5526
rect 6220 5516 6306 5526
rect 6014 5510 6306 5516
rect 6014 5476 6256 5510
rect 6290 5476 6306 5510
rect 6014 5468 6306 5476
rect 6014 5462 6098 5468
rect 6220 5462 6306 5468
rect 5946 5260 5986 5340
rect 6872 5268 6940 5280
rect 6872 5260 6888 5268
rect 5946 5248 6888 5260
rect 5946 5220 6458 5248
rect 6440 5214 6458 5220
rect 6492 5234 6888 5248
rect 6922 5234 6940 5268
rect 6492 5220 6940 5234
rect 6492 5214 6510 5220
rect 6440 5200 6510 5214
rect 5952 4930 6408 4946
rect 5952 4906 6354 4930
rect 5952 4820 5992 4906
rect 6338 4896 6354 4906
rect 6388 4896 6408 4930
rect 6338 4882 6408 4896
rect 6018 4716 6102 4726
rect 6224 4716 6306 4726
rect 6018 4710 6306 4716
rect 6018 4676 6254 4710
rect 6288 4676 6306 4710
rect 6018 4668 6306 4676
rect 6018 4662 6102 4668
rect 6224 4662 6306 4668
rect 5950 4478 5990 4540
rect 5950 4438 6674 4478
rect 5950 4106 6600 4146
rect 5950 4042 5990 4106
rect 6018 3916 6102 3922
rect 6224 3916 6306 3922
rect 6018 3906 6306 3916
rect 6018 3872 6254 3906
rect 6288 3872 6306 3906
rect 6018 3866 6306 3872
rect 6018 3856 6102 3866
rect 6224 3856 6306 3866
rect 5950 3664 5990 3740
rect 5950 3624 6526 3664
rect 5950 3306 6452 3346
rect 5950 3242 5990 3306
rect 6018 3116 6102 3122
rect 6224 3116 6306 3122
rect 6018 3110 6306 3116
rect 6018 3076 6254 3110
rect 6288 3076 6306 3110
rect 6018 3066 6306 3076
rect 6018 3064 6102 3066
rect 6224 3064 6306 3066
rect 2978 3012 3030 3024
rect 2978 2978 2986 3012
rect 3020 2978 3030 3012
rect 2978 2966 3030 2978
rect 2980 1440 3022 2966
rect 5950 2786 5990 2940
rect 6336 2786 6378 2792
rect 5950 2780 6378 2786
rect 5950 2746 6342 2780
rect 6376 2746 6378 2780
rect 5950 2496 6378 2536
rect 5950 2442 5990 2496
rect 6018 2316 6102 2324
rect 6224 2316 6306 2324
rect 6018 2310 6306 2316
rect 6018 2272 6254 2310
rect 6288 2272 6306 2310
rect 6018 2266 6306 2272
rect 6018 2262 6102 2266
rect 6224 2262 6306 2266
rect 5950 1664 5990 2140
rect 6340 1882 6378 2496
rect 6412 2302 6452 3306
rect 6486 2524 6526 3624
rect 6560 2734 6600 4106
rect 6634 2946 6674 4438
rect 6634 2926 6684 2946
rect 6634 2892 6642 2926
rect 6676 2892 6684 2926
rect 6634 2878 6684 2892
rect 6560 2716 6622 2734
rect 6560 2682 6572 2716
rect 6610 2682 6622 2716
rect 6560 2666 6622 2682
rect 6486 2508 6550 2524
rect 6486 2474 6498 2508
rect 6536 2474 6550 2508
rect 6486 2456 6550 2474
rect 6412 2282 6476 2302
rect 6412 2248 6428 2282
rect 6466 2248 6476 2282
rect 6412 2234 6476 2248
rect 6340 1862 6388 1882
rect 6340 1828 6346 1862
rect 6380 1828 6388 1862
rect 6340 1814 6388 1828
rect 5949 1650 6015 1664
rect 5949 1616 5964 1650
rect 5998 1616 6015 1650
rect 5949 1598 6015 1616
rect 2980 1386 3114 1440
rect 3960 1376 4012 1392
rect 3958 1340 4012 1376
rect 3960 1260 4012 1340
rect 2834 1208 4012 1260
rect 4804 1166 4860 1378
rect 2744 1110 4860 1166
rect 2660 1024 3034 1072
rect 2986 682 3034 1024
rect 2986 634 3132 682
rect 2907 554 3061 571
rect 2907 520 3010 554
rect 3044 520 3061 554
rect 2907 505 3061 520
rect 2907 205 2973 505
rect 7544 205 7610 1316
rect 7671 986 7737 10522
rect 7671 952 7686 986
rect 7724 952 7737 986
rect 7671 941 7737 952
rect 2907 139 7610 205
<< viali >>
rect 2456 9640 2490 9674
rect 2552 6974 2586 7008
rect 5952 10190 5986 10228
rect 6366 9972 6404 10006
rect 6256 9472 6290 9510
rect 6440 9766 6478 9800
rect 6522 9550 6560 9584
rect 6254 8672 6288 8706
rect 6606 9330 6644 9364
rect 2654 4310 2688 4344
rect 2756 8306 2790 8340
rect 2664 1646 2698 1680
rect 6678 9118 6716 9152
rect 6254 7874 6288 7908
rect 6464 7320 6498 7358
rect 6254 7074 6288 7108
rect 6586 6836 6620 6870
rect 6686 6506 6720 6540
rect 6256 6276 6290 6310
rect 6576 6036 6610 6070
rect 6786 5730 6820 5764
rect 2842 5644 2876 5678
rect 6256 5476 6290 5510
rect 6458 5214 6492 5248
rect 6888 5234 6922 5268
rect 6354 4896 6388 4930
rect 6254 4676 6288 4710
rect 6254 3872 6288 3906
rect 6254 3076 6288 3110
rect 2986 2978 3020 3012
rect 6342 2746 6376 2780
rect 6254 2272 6288 2310
rect 6642 2892 6676 2926
rect 6572 2682 6610 2716
rect 6498 2474 6536 2508
rect 6428 2248 6466 2282
rect 6346 1828 6380 1862
rect 5964 1616 5998 1650
rect 3588 738 3622 772
rect 4461 738 4495 772
rect 3255 642 3289 676
rect 3985 638 4019 672
rect 4127 638 4161 672
rect 3010 520 3044 554
rect 7686 952 7724 986
<< metal1 >>
rect 5370 10758 7084 10760
rect 2249 10676 7084 10758
rect 2249 10659 5391 10676
rect 3654 10548 3692 10659
rect 3850 10511 4133 10549
rect 4502 10548 4540 10659
rect 5346 10550 5384 10659
rect 5703 10574 6748 10646
rect 5703 10550 5766 10574
rect 2420 10088 2656 10092
rect 2648 10000 2656 10088
rect 2556 9974 2656 10000
rect 4095 9974 4133 10511
rect 4698 10510 4947 10548
rect 4909 9974 4947 10510
rect 5542 10509 5766 10550
rect 5725 9974 5766 10509
rect 5940 10240 5992 10242
rect 5940 10228 6876 10240
rect 5940 10190 5952 10228
rect 5986 10190 6876 10228
rect 5940 10174 6876 10190
rect 5940 10172 5992 10174
rect 6356 10006 6876 10024
rect 6238 9974 6306 9976
rect 2556 9890 6306 9974
rect 6356 9972 6366 10006
rect 6404 9972 6876 10006
rect 6356 9956 6876 9972
rect 3064 9830 3108 9890
rect 3064 9814 3140 9830
rect 3064 9778 3108 9814
rect 2446 9682 2500 9686
rect 2402 9674 2500 9682
rect 2402 9640 2456 9674
rect 2490 9640 2500 9674
rect 2402 9630 2500 9640
rect 2446 9628 2500 9630
rect 2426 9480 3068 9524
rect 6238 9510 6306 9890
rect 6432 9800 6950 9818
rect 6432 9766 6440 9800
rect 6478 9766 6950 9800
rect 6432 9748 6950 9766
rect 6515 9584 6950 9604
rect 6515 9550 6522 9584
rect 6560 9550 6950 9584
rect 6515 9534 6950 9550
rect 2426 9426 2526 9480
rect 2392 9424 2526 9426
rect 2426 9418 2526 9424
rect 6238 9472 6256 9510
rect 6290 9472 6306 9510
rect 2556 9220 3116 9228
rect 2556 9138 2564 9220
rect 2644 9176 3148 9220
rect 2644 9138 2654 9176
rect 2556 9130 2654 9138
rect 3064 9030 3108 9176
rect 3064 8986 3136 9030
rect 3064 8978 3108 8986
rect 2956 8672 3066 8734
rect 6238 8706 6306 9472
rect 6599 9364 6950 9384
rect 6599 9330 6606 9364
rect 6644 9330 6950 9364
rect 6599 9314 6950 9330
rect 6672 9152 6950 9172
rect 6672 9118 6678 9152
rect 6716 9118 6950 9152
rect 6672 9104 6950 9118
rect 6238 8672 6254 8706
rect 6288 8672 6306 8706
rect 2956 8628 3023 8672
rect 2426 8614 3023 8628
rect 2426 8560 2448 8614
rect 2502 8570 3023 8614
rect 2502 8560 2526 8570
rect 2426 8550 2526 8560
rect 2554 8464 2654 8480
rect 2554 8410 2572 8464
rect 2626 8446 2654 8464
rect 2626 8410 3190 8446
rect 2554 8394 3190 8410
rect 3064 8386 3108 8394
rect 3064 8376 3140 8386
rect 2740 8350 2800 8352
rect 2422 8340 2800 8350
rect 2422 8306 2756 8340
rect 2790 8306 2800 8340
rect 2422 8298 2800 8306
rect 2740 8294 2800 8298
rect 3064 8230 3108 8376
rect 3064 8220 3134 8230
rect 3064 8178 3108 8220
rect 2426 7934 2526 7996
rect 2426 7872 3068 7934
rect 6238 7908 6306 8672
rect 6238 7874 6254 7908
rect 6288 7874 6306 7908
rect 3064 7564 3136 7590
rect 3064 7442 3126 7564
rect 3064 7428 3136 7442
rect 2434 7420 3136 7428
rect 2434 7406 3088 7420
rect 2434 7394 3190 7406
rect 2642 7374 3190 7394
rect 2426 7134 2526 7150
rect 2426 7126 3068 7134
rect 2426 7074 2446 7126
rect 2500 7074 3068 7126
rect 2426 7072 3068 7074
rect 6238 7108 6306 7874
rect 6448 8892 6896 8960
rect 6448 7358 6516 8892
rect 6448 7320 6464 7358
rect 6498 7320 6516 7358
rect 6448 7312 6516 7320
rect 6570 8678 6894 8746
rect 6238 7074 6254 7108
rect 6288 7074 6306 7108
rect 2426 7050 2526 7072
rect 2442 7008 2598 7018
rect 2442 6974 2552 7008
rect 2586 6974 2598 7008
rect 2442 6966 2598 6974
rect 3064 6790 3116 6828
rect 3064 6776 3136 6790
rect 3064 6630 3116 6776
rect 2556 6622 3136 6630
rect 2556 6540 2564 6622
rect 2644 6616 3136 6622
rect 2644 6578 3116 6616
rect 2644 6540 2654 6578
rect 2556 6532 2654 6540
rect 3011 6333 3068 6334
rect 2426 6240 2526 6254
rect 3011 6240 3069 6333
rect 2426 6236 3069 6240
rect 2426 6184 2448 6236
rect 2504 6184 3069 6236
rect 2426 6182 3069 6184
rect 6238 6310 6306 7074
rect 6570 6870 6638 8678
rect 6570 6836 6586 6870
rect 6620 6836 6638 6870
rect 6570 6824 6638 6836
rect 6668 8476 6896 8544
rect 6238 6276 6256 6310
rect 6290 6276 6306 6310
rect 2426 6166 2526 6182
rect 2629 6014 3122 6028
rect 2556 5970 3190 6014
rect 3064 5778 3108 5970
rect 2834 5686 2888 5690
rect 2438 5678 2888 5686
rect 2438 5644 2842 5678
rect 2876 5644 2888 5678
rect 2438 5634 2888 5644
rect 2834 5632 2888 5634
rect 2425 5482 3064 5524
rect 6238 5510 6306 6276
rect 6668 6540 6736 8476
rect 6668 6506 6686 6540
rect 6720 6506 6736 6540
rect 2426 5430 2526 5482
rect 2394 5428 2526 5430
rect 2426 5328 2526 5428
rect 6238 5476 6256 5510
rect 6290 5476 6306 5510
rect 2556 5224 3108 5228
rect 2556 5142 2562 5224
rect 2642 5184 3108 5224
rect 2642 5142 2654 5184
rect 2556 5140 2654 5142
rect 3064 4978 3108 5184
rect 2426 4616 2526 4630
rect 2426 4562 2446 4616
rect 2500 4612 2526 4616
rect 3054 4612 3094 4724
rect 2500 4572 3094 4612
rect 6238 4710 6306 5476
rect 6558 6070 6628 6084
rect 6558 6036 6576 6070
rect 6610 6036 6628 6070
rect 6440 5248 6510 5260
rect 6440 5214 6458 5248
rect 6492 5214 6510 5248
rect 6238 4676 6254 4710
rect 6288 4676 6306 4710
rect 2500 4562 2526 4572
rect 2426 4548 2526 4562
rect 2416 4344 2704 4354
rect 2416 4310 2654 4344
rect 2688 4310 2704 4344
rect 2416 4302 2704 4310
rect 3064 4220 3108 4428
rect 2556 4214 3108 4220
rect 2556 4132 2564 4214
rect 2644 4176 3108 4214
rect 2644 4132 2654 4176
rect 2556 4126 2654 4132
rect 2485 4009 2527 4093
rect 2459 4007 2527 4009
rect 2425 3924 2527 4007
rect 2425 3882 3072 3924
rect 6238 3906 6306 4676
rect 6238 3872 6254 3906
rect 6288 3872 6306 3906
rect 3064 3432 3108 3628
rect 2336 3378 3108 3432
rect 2336 3332 2654 3378
rect 2427 3152 2525 3169
rect 2427 3098 2448 3152
rect 2502 3124 2525 3152
rect 2502 3098 3066 3124
rect 2427 3082 3066 3098
rect 6238 3110 6306 3872
rect 6238 3076 6254 3110
rect 6288 3076 6306 3110
rect 6338 4930 6408 4944
rect 6338 4896 6354 4930
rect 6388 4896 6408 4930
rect 6338 3161 6408 4896
rect 6440 3361 6510 5214
rect 6558 3573 6628 6036
rect 6668 3786 6736 6506
rect 6768 8286 6896 8334
rect 6768 8266 6950 8286
rect 6768 5764 6836 8266
rect 6768 5730 6786 5764
rect 6820 5730 6836 5764
rect 6768 5716 6836 5730
rect 6872 8068 6896 8076
rect 6872 5268 6940 8068
rect 6872 5234 6888 5268
rect 6922 5234 6940 5268
rect 6872 5220 6940 5234
rect 6668 3718 6930 3786
rect 6558 3503 6931 3573
rect 6440 3291 6931 3361
rect 6338 3091 6931 3161
rect 2978 3022 3030 3024
rect 2442 3012 3030 3022
rect 2442 2978 2986 3012
rect 3020 2978 3030 3012
rect 2442 2970 3030 2978
rect 2978 2966 3030 2970
rect 2556 2754 2656 2764
rect 2556 2672 2566 2754
rect 2646 2740 2656 2754
rect 3064 2740 3108 2824
rect 2646 2696 3108 2740
rect 2646 2672 2656 2696
rect 2556 2664 2656 2672
rect 3064 2578 3108 2696
rect 2426 2254 2526 2262
rect 2426 2172 2436 2254
rect 2516 2236 2526 2254
rect 3060 2236 3104 2324
rect 6238 2310 6306 3076
rect 6634 2926 6930 2946
rect 6634 2892 6642 2926
rect 6676 2892 6930 2926
rect 6634 2878 6930 2892
rect 6238 2272 6254 2310
rect 6288 2272 6306 2310
rect 6238 2262 6306 2272
rect 6336 2780 6390 2792
rect 6336 2746 6342 2780
rect 6376 2746 6390 2780
rect 2516 2192 3104 2236
rect 2516 2172 2526 2192
rect 2426 2162 2526 2172
rect 2336 2028 2656 2100
rect 6336 2088 6390 2746
rect 6560 2716 6930 2734
rect 6560 2682 6572 2716
rect 6610 2682 6930 2716
rect 6560 2666 6930 2682
rect 6486 2508 6930 2524
rect 6486 2474 6498 2508
rect 6536 2474 6930 2508
rect 6486 2456 6930 2474
rect 6418 2282 6932 2302
rect 6418 2248 6428 2282
rect 6466 2248 6932 2282
rect 6418 2234 6932 2248
rect 6336 2087 6922 2088
rect 6336 2033 6927 2087
rect 6336 2028 6922 2033
rect 2336 2000 3120 2028
rect 6336 2020 6930 2028
rect 2556 1984 3120 2000
rect 2556 1888 2656 1984
rect 2556 1788 5345 1888
rect 6340 1862 6930 1882
rect 6340 1828 6346 1862
rect 6380 1828 6930 1862
rect 6340 1814 6930 1828
rect 2660 1690 2710 1692
rect 2418 1680 2710 1690
rect 2418 1646 2664 1680
rect 2698 1646 2710 1680
rect 2418 1638 2710 1646
rect 2660 1634 2710 1638
rect 2390 1428 2526 1434
rect 2424 1424 2526 1428
rect 2426 1234 2526 1332
rect 3635 1309 3673 1788
rect 3428 1271 3673 1309
rect 4489 1308 4527 1788
rect 3232 1234 3270 1268
rect 4080 1234 4118 1272
rect 4276 1270 4527 1308
rect 4915 1234 4969 1357
rect 5307 1312 5345 1788
rect 5949 1650 6862 1664
rect 5949 1616 5964 1650
rect 5998 1616 6862 1650
rect 5949 1598 6862 1616
rect 5120 1274 5345 1312
rect 2426 1166 4969 1234
rect 5287 1264 5345 1274
rect 5287 1192 6796 1264
rect 3072 1062 4618 1166
rect 4915 1130 4969 1166
rect 6970 1130 6994 1144
rect 4915 1076 7032 1130
rect 2389 968 2889 1027
rect 3742 984 4618 1062
rect 5467 986 7739 996
rect 2830 912 2889 968
rect 5467 952 7686 986
rect 7724 952 7739 986
rect 5467 942 7739 952
rect 5467 919 5521 942
rect 2830 853 4035 912
rect 3574 772 3798 780
rect 3574 738 3588 772
rect 3622 738 3798 772
rect 3574 728 3798 738
rect 3240 676 3308 686
rect 3240 642 3255 676
rect 3289 642 3308 676
rect 3240 620 3308 642
rect 3241 572 3307 620
rect 2995 554 3307 572
rect 2995 520 3010 554
rect 3044 520 3307 554
rect 2995 506 3307 520
rect 3746 546 3798 728
rect 3976 672 4035 853
rect 3976 638 3985 672
rect 4019 638 4035 672
rect 3976 623 4035 638
rect 4111 865 5521 919
rect 4111 678 4165 865
rect 4448 772 7746 782
rect 4448 738 4461 772
rect 4495 738 7746 772
rect 4448 730 7746 738
rect 4111 672 4168 678
rect 4111 638 4127 672
rect 4161 638 4168 672
rect 4111 630 4168 638
rect 4111 617 4165 630
rect 2995 505 3061 506
rect 3746 494 7750 546
rect 2557 392 3104 416
rect 2557 346 2574 392
rect 2556 338 2574 346
rect 2628 384 3104 392
rect 2628 350 3103 384
rect 3718 350 4617 416
rect 2628 346 3104 350
rect 3702 346 4617 350
rect 2628 338 4617 346
rect 2556 314 4617 338
<< via1 >>
rect 2564 9138 2644 9220
rect 2448 8560 2502 8614
rect 2572 8410 2626 8464
rect 2446 7074 2500 7126
rect 2564 6540 2644 6622
rect 2448 6184 2504 6236
rect 2562 5142 2642 5224
rect 2446 4562 2500 4616
rect 2564 4132 2644 4214
rect 2448 3098 2502 3152
rect 2566 2672 2646 2754
rect 2436 2172 2516 2254
rect 2574 338 2628 392
<< metal2 >>
rect 213 10760 273 10764
rect 12 10660 56 10760
rect 102 10670 146 10760
rect 2426 10752 2526 10766
rect 2556 10748 2654 10766
rect 2556 392 2654 865
rect 2556 338 2574 392
rect 2628 338 2654 392
rect 2556 317 2654 338
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 3072 0 1 367
box -38 -49 710 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_1
timestamp 1626515395
transform 1 0 3944 0 1 363
box -38 -49 710 715
use ROM_cell  ROM_cell_1
timestamp 1641148104
transform 1 0 7246 0 -1 2112
box -522 -1846 364 1036
use ROM_cell  ROM_cell_0
timestamp 1641148104
transform 1 0 7266 0 1 9726
box -522 -1846 364 1036
use sparse_decoder  sparse_decoder_0
timestamp 1641072977
transform 1 0 3064 0 1 9472
box -176 -8374 3128 1288
use asyn_rst_8_gray_counter  asyn_rst_8_gray_counter_0
timestamp 1640932070
transform 1 0 174 0 1 9324
box -174 -9324 2481 1438
<< labels >>
rlabel metal2 30 10760 30 10760 1 clk
port 3 n
rlabel metal2 122 10760 122 10760 1 RST_bar
port 4 n
rlabel metal2 242 10764 242 10764 1 EN
port 5 n
rlabel metal2 2474 10766 2474 10766 1 VDD
port 7 n
rlabel metal2 2604 10766 2604 10766 1 GND
port 6 n
rlabel metal1 7746 756 7746 756 3 sine_out
port 1 e
rlabel metal1 7750 520 7750 520 3 cos_out
port 2 e
<< end >>
