* NGSPICE file created from user_proj.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

.subckt user_proj io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i vccd1 vssd1
+ vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vssa2_uq0 vssa2_uq1 vssa2_uq2 vssa2_uq3 vssa2_uq4
+ vssa1_uq0 vssa1_uq1 vssa1_uq2 vssa1_uq3 vssa1_uq4 vssd2_uq0 vssd2_uq1 vssd2_uq2
+ vssd2_uq3 vssd2_uq4 vdda2_uq0 vdda2_uq1 vdda2_uq2 vdda2_uq3 vdda2_uq4 vdda1_uq0
+ vdda1_uq1 vdda1_uq2 vdda1_uq3 vdda1_uq4 vccd2_uq0 vccd2_uq1 vccd2_uq2 vccd2_uq3
+ vccd2_uq4
XFILLER_100_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09671_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09671_/Y sky130_fd_sc_hd__inv_2
X_06883_ _06958_/A vssd1 vssd1 vccd1 vccd1 _06883_/X sky130_fd_sc_hd__buf_1
XFILLER_94_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08622_ _13763_/Q _08618_/X _08530_/X _08619_/X _08620_/X vssd1 vssd1 vccd1 vccd1
+ _13763_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ _08957_/A vssd1 vssd1 vccd1 vccd1 _08553_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07504_ _14319_/Q _07499_/X _07327_/X _07501_/X _07503_/X vssd1 vssd1 vccd1 vccd1
+ _14319_/D sky130_fd_sc_hd__o221a_1
X_08484_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08565_/A sky130_fd_sc_hd__inv_2
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07435_ _14354_/Q _07432_/X _07336_/X _07433_/X _07434_/X vssd1 vssd1 vccd1 vccd1
+ _14354_/D sky130_fd_sc_hd__o221a_1
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07366_ _14382_/Q _07361_/X _07365_/X _07363_/X _07359_/X vssd1 vssd1 vccd1 vccd1
+ _14382_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09105_ _13518_/Q _09103_/X _08945_/X _09104_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _13518_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07297_ _14408_/Q _07290_/X _06837_/X _07291_/X _07295_/X vssd1 vssd1 vccd1 vccd1
+ _14408_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _09036_/A vssd1 vssd1 vccd1 vccd1 _09036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _09901_/A _09901_/B _09937_/Y vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ _13299_/Q vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__inv_2
XFILLER_150_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11900_ _13932_/Q vssd1 vssd1 vccd1 vccd1 _11900_/Y sky130_fd_sc_hd__inv_2
XPHY_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12531_/X input339/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _12236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11831_ _11831_/A vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14550_ _14629_/CLK _14550_/D vssd1 vssd1 vccd1 vccd1 _14550_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11762_ _13727_/Q _11642_/X _14046_/Q _11663_/X _11761_/X vssd1 vssd1 vccd1 vccd1
+ _11762_/X sky130_fd_sc_hd__a221o_4
XPHY_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13501_ _14094_/CLK _13501_/D vssd1 vssd1 vccd1 vccd1 _13501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10713_ _13985_/Q vssd1 vssd1 vccd1 vccd1 _10713_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14481_/CLK _14481_/D vssd1 vssd1 vccd1 vccd1 _14481_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11693_/A vssd1 vssd1 vccd1 vccd1 _11693_/X sky130_fd_sc_hd__buf_2
XPHY_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _14143_/CLK _13432_/D vssd1 vssd1 vccd1 vccd1 _13432_/Q sky130_fd_sc_hd__dfxtp_1
X_10644_ _10644_/A _10644_/B _10644_/C _10644_/D vssd1 vssd1 vccd1 vccd1 _10644_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10575_ _13826_/Q vssd1 vssd1 vccd1 vccd1 _10575_/Y sky130_fd_sc_hd__inv_2
X_13363_ _14639_/CLK _13363_/D vssd1 vssd1 vccd1 vccd1 _13363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12314_ _10644_/Y _14529_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _13877_/CLK _13294_/D vssd1 vssd1 vccd1 vccd1 _13294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12176_ vssd1 vssd1 vccd1 vccd1 _12176_/HI _12176_/LO sky130_fd_sc_hd__conb_1
XFILLER_170_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ _13955_/Q vssd1 vssd1 vccd1 vccd1 _11127_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11058_ _14499_/Q vssd1 vssd1 vccd1 vccd1 _11058_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10009_ _13375_/Q _10008_/B _10010_/A vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07220_ _14450_/Q _07217_/X _07073_/X _07218_/X _07213_/X vssd1 vssd1 vccd1 vccd1
+ _14450_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07151_ _14486_/Q _07144_/X _06837_/X _07145_/X _07147_/X vssd1 vssd1 vccd1 vccd1
+ _14486_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ _14522_/Q _07014_/A _06850_/B _07017_/A _07079_/X vssd1 vssd1 vccd1 vccd1
+ _14522_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput401 _12201_/X vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput412 _12091_/LO vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput423 _12239_/A vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput434 _12249_/A vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput445 _12097_/LO vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput456 _12243_/X vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput467 _10126_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput478 _12111_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput489 _12121_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07984_ _14076_/Q _07982_/X _07746_/X _07983_/X _07978_/X vssd1 vssd1 vccd1 vccd1
+ _14076_/D sky130_fd_sc_hd__o221a_1
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ _09701_/A _09722_/X _09701_/A _09722_/X vssd1 vssd1 vccd1 vccd1 _09723_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06935_ _06935_/A _06935_/B vssd1 vssd1 vccd1 vccd1 _14579_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09654_ _09613_/X _09653_/Y _09613_/X _09653_/Y vssd1 vssd1 vccd1 vccd1 _09654_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06866_ _06857_/X _12285_/X _06865_/X _06861_/X vssd1 vssd1 vccd1 vccd1 _06867_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ _13773_/Q _08599_/X _08505_/X _08601_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _13773_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09585_ _09583_/X _09582_/X _13261_/Q _09584_/X vssd1 vssd1 vccd1 vccd1 _13229_/D
+ sky130_fd_sc_hd__o22a_1
X_06797_ _14615_/Q _06787_/X _06796_/X _06790_/X _06785_/X vssd1 vssd1 vccd1 vccd1
+ _14615_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08536_ _08942_/A vssd1 vssd1 vccd1 vccd1 _08536_/X sky130_fd_sc_hd__clkbuf_4
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _13828_/Q _08460_/X _08171_/X _08461_/X _08465_/X vssd1 vssd1 vccd1 vccd1
+ _13828_/D sky130_fd_sc_hd__o221a_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ _14362_/Q _07411_/X _07313_/X _07414_/X _07415_/X vssd1 vssd1 vccd1 vccd1
+ _14362_/D sky130_fd_sc_hd__o221a_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08398_ _13866_/Q _08396_/X _08175_/X _08397_/X _08392_/X vssd1 vssd1 vccd1 vccd1
+ _13866_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07349_ _08137_/A vssd1 vssd1 vccd1 vccd1 _07349_/X sky130_fd_sc_hd__buf_2
XFILLER_136_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _13542_/Q _10206_/X _13783_/Q _10209_/X vssd1 vssd1 vccd1 vccd1 _10360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _09036_/A vssd1 vssd1 vccd1 vccd1 _09019_/X sky130_fd_sc_hd__buf_2
X_10291_ _13898_/Q vssd1 vssd1 vccd1 vccd1 _10291_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12030_ _12030_/A _12030_/B _12030_/C _12030_/D vssd1 vssd1 vccd1 vccd1 _12030_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _14100_/CLK _13981_/D vssd1 vssd1 vccd1 vccd1 _13981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ _12547_/X input357/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12526_/X _12862_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14637_/CLK _14602_/D vssd1 vssd1 vccd1 vccd1 _14602_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11812_/Y _11683_/X _11813_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11814_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12794_ _09537_/X _12793_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12794_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14611_/CLK _14533_/D vssd1 vssd1 vccd1 vccd1 _14533_/Q sky130_fd_sc_hd__dfxtp_1
X_11745_ _11743_/Y _11637_/X _11744_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _11745_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464_ _14595_/CLK _14464_/D vssd1 vssd1 vccd1 vccd1 _14464_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11672_/Y _11673_/X _11674_/Y _11675_/X vssd1 vssd1 vccd1 vccd1 _11676_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13415_ _14178_/CLK _13415_/D vssd1 vssd1 vccd1 vccd1 _13415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10627_ _14607_/Q vssd1 vssd1 vccd1 vccd1 _10627_/Y sky130_fd_sc_hd__inv_2
X_14395_ _14629_/CLK _14395_/D vssd1 vssd1 vccd1 vccd1 _14395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13346_ _14538_/CLK _13346_/D vssd1 vssd1 vccd1 vccd1 _13346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10558_ _10556_/Y _10512_/X _10557_/Y _10515_/X vssd1 vssd1 vccd1 vccd1 _10558_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_196_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13277_ _14573_/CLK _13277_/D vssd1 vssd1 vccd1 vccd1 _13277_/Q sky130_fd_sc_hd__dfxtp_4
X_10489_ _10476_/Y _10478_/X _10479_/Y _10481_/X _10488_/X vssd1 vssd1 vccd1 vccd1
+ _10518_/B sky130_fd_sc_hd__o221a_2
XFILLER_100_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12228_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12159_ vssd1 vssd1 vccd1 vccd1 _12159_/HI _12159_/LO sky130_fd_sc_hd__conb_1
XFILLER_25_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06720_ _14635_/Q _06530_/X _06719_/X _06716_/X _06723_/C1 vssd1 vssd1 vccd1 vccd1
+ _14635_/D sky130_fd_sc_hd__o221a_1
XFILLER_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06651_ _06829_/B vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__inv_2
XFILLER_209_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09370_ _09370_/A _12799_/X vssd1 vssd1 vccd1 vccd1 _13358_/D sky130_fd_sc_hd__and2_1
X_06582_ _06609_/A vssd1 vssd1 vccd1 vccd1 _06582_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08321_ _08329_/A vssd1 vssd1 vccd1 vccd1 _08321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08252_ _13947_/Q _08246_/X _08167_/X _08247_/X _08249_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07203_ _14461_/Q _07201_/X _06789_/X _07202_/X _07197_/X vssd1 vssd1 vccd1 vccd1
+ _14461_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _08183_/A vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__buf_4
XFILLER_203_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07134_ _14497_/Q _07127_/X _07058_/X _07128_/X _07131_/X vssd1 vssd1 vccd1 vccd1
+ _14497_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07065_ _14533_/Q _07061_/X _06810_/X _07062_/X _07063_/X vssd1 vssd1 vccd1 vccd1
+ _14533_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07967_ _08000_/A vssd1 vssd1 vccd1 vccd1 _07967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _06902_/Y _14584_/Q _14588_/Q _06915_/Y vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_5_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06918_ _06918_/A vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ _14124_/Q _07892_/X _07723_/X _07894_/X _07897_/X vssd1 vssd1 vccd1 vccd1
+ _14124_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09637_ _09637_/A vssd1 vssd1 vccd1 vccd1 _09637_/Y sky130_fd_sc_hd__inv_2
X_06849_ _08985_/A vssd1 vssd1 vccd1 vccd1 _06850_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_99_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09568_ _09557_/X _09567_/X _13267_/Q _09558_/X vssd1 vssd1 vccd1 vccd1 _13235_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _08922_/A vssd1 vssd1 vccd1 vccd1 _08519_/X sky130_fd_sc_hd__clkbuf_4
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _13262_/Q _09493_/X _12257_/X _09494_/X vssd1 vssd1 vccd1 vccd1 _13262_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11530_ _14509_/Q vssd1 vssd1 vccd1 vccd1 _11530_/Y sky130_fd_sc_hd__inv_2
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ _11461_/A vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13200_ _13368_/CLK _13200_/D vssd1 vssd1 vccd1 vccd1 _13200_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ _14252_/Q vssd1 vssd1 vccd1 vccd1 _10412_/Y sky130_fd_sc_hd__inv_2
X_14180_ _14183_/CLK _14180_/D vssd1 vssd1 vccd1 vccd1 _14180_/Q sky130_fd_sc_hd__dfxtp_1
X_11392_ _11390_/Y _11223_/X _11391_/Y _11225_/X vssd1 vssd1 vccd1 vccd1 _11392_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _12643_/X _13130_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _13659_/Q vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10274_ _10264_/Y _10178_/X _10267_/X _10270_/X _10273_/X vssd1 vssd1 vccd1 vccd1
+ _10298_/C sky130_fd_sc_hd__o2111a_4
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13062_ _13061_/X _12610_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _14637_/Q vssd1 vssd1 vccd1 vccd1 _12013_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13964_ _14110_/CLK _13964_/D vssd1 vssd1 vccd1 vccd1 _13964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12915_ _12539_/X _12914_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12915_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13895_ _14130_/CLK _13895_/D vssd1 vssd1 vccd1 vccd1 _13895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12846_ _12522_/X _12845_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12846_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12777_ _09524_/X _12776_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14516_ _14637_/CLK _14516_/D vssd1 vssd1 vccd1 vccd1 _14516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _13609_/Q vssd1 vssd1 vccd1 vccd1 _11728_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14447_ _14481_/CLK _14447_/D vssd1 vssd1 vccd1 vccd1 _14447_/Q sky130_fd_sc_hd__dfxtp_1
X_11659_ _13530_/Q vssd1 vssd1 vccd1 vccd1 _11659_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14378_ _14627_/CLK _14378_/D vssd1 vssd1 vccd1 vccd1 _14378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13329_ _14639_/CLK _13329_/D vssd1 vssd1 vccd1 vccd1 _13329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08870_ _13630_/Q _08868_/X _08553_/X _08869_/X _08863_/X vssd1 vssd1 vccd1 vccd1
+ _13630_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07821_ _07856_/A vssd1 vssd1 vccd1 vccd1 _07821_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater701 _13085_/S vssd1 vssd1 vccd1 vccd1 _13145_/S sky130_fd_sc_hd__buf_8
XFILLER_6_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07752_ _14191_/Q _07745_/X _07751_/X _07747_/X _07743_/X vssd1 vssd1 vccd1 vccd1
+ _14191_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06703_ _12396_/S _09035_/A vssd1 vssd1 vccd1 vccd1 _06703_/X sky130_fd_sc_hd__and2_1
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07683_ _14220_/Q _07679_/X _07379_/X _07680_/X _07676_/X vssd1 vssd1 vccd1 vccd1
+ _14220_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09422_ _09426_/A _13027_/X vssd1 vssd1 vccd1 vccd1 _13317_/D sky130_fd_sc_hd__and2_1
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06634_ _06573_/X _06633_/X _06573_/A _06633_/X vssd1 vssd1 vccd1 vccd1 _06634_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_168_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ _09357_/A _12871_/X vssd1 vssd1 vccd1 vccd1 _13372_/D sky130_fd_sc_hd__and2_1
X_06565_ _06565_/A vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08304_ _13920_/Q _08302_/X _08137_/X _08303_/X _08297_/X vssd1 vssd1 vccd1 vccd1
+ _13920_/D sky130_fd_sc_hd__o221a_1
XFILLER_166_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _09326_/A vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__clkbuf_4
X_06496_ _06496_/A vssd1 vssd1 vccd1 vccd1 _06497_/B sky130_fd_sc_hd__inv_2
XFILLER_178_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08235_ _13956_/Q _08229_/X _08144_/X _08230_/X _08231_/X vssd1 vssd1 vccd1 vccd1
+ _13956_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08166_ _13987_/Q _08161_/X _08165_/X _08163_/X _08159_/X vssd1 vssd1 vccd1 vccd1
+ _13987_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07117_ _14507_/Q _07111_/X _06763_/X _07112_/X _07114_/X vssd1 vssd1 vccd1 vccd1
+ _14507_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08097_ _08097_/A vssd1 vssd1 vccd1 vccd1 _08097_/X sky130_fd_sc_hd__buf_2
XFILLER_146_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07048_ _14543_/Q _07044_/X _06775_/X _07045_/X _07046_/X vssd1 vssd1 vccd1 vccd1
+ _14543_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _09138_/A vssd1 vssd1 vccd1 vccd1 _09036_/A sky130_fd_sc_hd__buf_2
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _13206_/Q _10775_/X _14029_/Q _10957_/X _10960_/X vssd1 vssd1 vccd1 vccd1
+ _10961_/X sky130_fd_sc_hd__a221o_4
XFILLER_99_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ _09560_/X input336/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13680_ _14143_/CLK _13680_/D vssd1 vssd1 vccd1 vccd1 _13680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10892_ _10890_/Y _10704_/X _10891_/Y _10706_/X vssd1 vssd1 vccd1 vccd1 _10892_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ _13329_/Q _12630_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12562_ _13300_/Q _12561_/X input39/X vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__mux2_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14301_ _14305_/CLK _14301_/D vssd1 vssd1 vccd1 vccd1 _14301_/Q sky130_fd_sc_hd__dfxtp_1
X_11513_ _11508_/Y _11397_/X _11509_/Y _11399_/X _11512_/X vssd1 vssd1 vccd1 vccd1
+ _11549_/A sky130_fd_sc_hd__o221a_2
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12492_/X _06975_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__mux2_2
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14232_ _14595_/CLK _14232_/D vssd1 vssd1 vccd1 vccd1 _14232_/Q sky130_fd_sc_hd__dfxtp_1
X_11444_ _14312_/Q vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14163_ _14291_/CLK _14163_/D vssd1 vssd1 vccd1 vccd1 _14163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11375_ _13215_/Q _11249_/X _14038_/Q _11193_/X _11374_/X vssd1 vssd1 vccd1 vccd1
+ _11375_/X sky130_fd_sc_hd__a221o_4
XFILLER_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _13113_/X _12635_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__mux2_1
X_10326_ _10321_/Y _10214_/X _10322_/Y _10217_/X _10325_/X vssd1 vssd1 vccd1 vccd1
+ _10339_/B sky130_fd_sc_hd__o221a_2
XFILLER_49_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14094_ _14094_/CLK _14094_/D vssd1 vssd1 vccd1 vccd1 _14094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13045_ _12602_/X _13044_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13045_/X sky130_fd_sc_hd__mux2_1
X_10257_ _13423_/Q vssd1 vssd1 vccd1 vccd1 _10257_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10188_ _10188_/A vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13947_ _14107_/CLK _13947_/D vssd1 vssd1 vccd1 vccd1 _13947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13878_ _13996_/CLK _13878_/D vssd1 vssd1 vccd1 vccd1 _13878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _12518_/X _12828_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08020_ _08813_/A vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__buf_2
XFILLER_11_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09971_ _09971_/A vssd1 vssd1 vccd1 vccd1 _09972_/B sky130_fd_sc_hd__inv_2
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ _08922_/A vssd1 vssd1 vccd1 vccd1 _08922_/X sky130_fd_sc_hd__buf_6
XFILLER_83_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08853_ _08869_/A vssd1 vssd1 vccd1 vccd1 _08853_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _08411_/A _07878_/B _08814_/C _08091_/D vssd1 vssd1 vccd1 vccd1 _11691_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_22_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _08793_/A vssd1 vssd1 vccd1 vccd1 _08784_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _14198_/Q _07732_/X _07733_/X _07734_/X _07730_/X vssd1 vssd1 vccd1 vccd1
+ _14198_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07666_/X sky130_fd_sc_hd__buf_2
XFILLER_80_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09405_ _09407_/A _13103_/X vssd1 vssd1 vccd1 vccd1 _13330_/D sky130_fd_sc_hd__and2_1
XFILLER_41_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06617_ input93/X vssd1 vssd1 vccd1 vccd1 _06617_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07597_ _07605_/A vssd1 vssd1 vccd1 vccd1 _07597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09336_ _09336_/A vssd1 vssd1 vccd1 vccd1 _09509_/A sky130_fd_sc_hd__buf_2
X_06548_ _06542_/X _06547_/X _06542_/X _06547_/X vssd1 vssd1 vccd1 vccd1 _06548_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09267_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09267_/X sky130_fd_sc_hd__buf_2
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08218_ _13967_/Q _08211_/X _08217_/X _08213_/X _08214_/X vssd1 vssd1 vccd1 vccd1
+ _13967_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09198_ _13463_/Q _09135_/A _08983_/X _09137_/A _09196_/X vssd1 vssd1 vccd1 vccd1
+ _13463_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08149_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11160_ _14073_/Q vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10111_ _10111_/A _12466_/X vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__nor2_8
XFILLER_161_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11091_ _14110_/Q vssd1 vssd1 vccd1 vccd1 _11091_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput301 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _06502_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ _13363_/Q _09984_/B _09985_/A vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__o21a_1
Xinput312 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _06495_/C sky130_fd_sc_hd__clkbuf_1
XPHY_7333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput323 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _06507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput334 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input334/X sky130_fd_sc_hd__clkbuf_4
XPHY_7355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput345 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 input345/X sky130_fd_sc_hd__buf_6
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput356 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input356/X sky130_fd_sc_hd__clkbuf_4
XPHY_7377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput367 wbs_we_i vssd1 vssd1 vccd1 vccd1 _12853_/S sky130_fd_sc_hd__buf_6
XFILLER_40_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _13996_/CLK _13801_/D vssd1 vssd1 vccd1 vccd1 _13801_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11993_ _13655_/Q vssd1 vssd1 vccd1 vccd1 _11993_/Y sky130_fd_sc_hd__inv_2
XPHY_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13732_ _14056_/CLK _13732_/D vssd1 vssd1 vccd1 vccd1 _13732_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _11416_/A vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13663_ _14047_/CLK _13663_/D vssd1 vssd1 vccd1 vccd1 _13663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10875_ _13474_/Q vssd1 vssd1 vccd1 vccd1 _10875_/Y sky130_fd_sc_hd__inv_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _13322_/Q _12613_/X input39/X vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__mux2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13594_ _14188_/CLK _13594_/D vssd1 vssd1 vccd1 vccd1 _13594_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12545_ _13293_/Q _12544_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12476_ _12509_/X _06957_/Y _12476_/S vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ _14291_/CLK _14215_/D vssd1 vssd1 vccd1 vccd1 _14215_/Q sky130_fd_sc_hd__dfxtp_1
X_11427_ _11423_/Y _11424_/X _11425_/Y _11426_/X vssd1 vssd1 vccd1 vccd1 _11427_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 _10993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _14146_/CLK _14146_/D vssd1 vssd1 vccd1 vccd1 _14146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11358_ _13641_/Q vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10309_ _13743_/Q vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14077_ _14305_/CLK _14077_/D vssd1 vssd1 vccd1 vccd1 _14077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _13522_/Q vssd1 vssd1 vccd1 vccd1 _11289_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13028_ _12594_/X input351/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13028_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07520_ _14309_/Q _07516_/X _07352_/X _07517_/X _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14309_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07451_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07382_ _14375_/Q _07373_/X _07381_/X _07375_/X _07371_/X vssd1 vssd1 vccd1 vccd1
+ _14375_/D sky130_fd_sc_hd__o221a_1
XFILLER_56_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09121_ _13508_/Q _09119_/X _08970_/X _09120_/X _09117_/X vssd1 vssd1 vccd1 vccd1
+ _13508_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _13546_/Q _09048_/X _09051_/X _09049_/X _09045_/X vssd1 vssd1 vccd1 vccd1
+ _13546_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08003_ _08017_/A vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _13302_/Q _09952_/Y _09897_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08905_ _08956_/A vssd1 vssd1 vccd1 vccd1 _08905_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09885_ _09885_/A _09958_/A vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__or2_1
XFILLER_150_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08836_ _13650_/Q _08832_/X _08833_/X _08835_/X _08823_/X vssd1 vssd1 vccd1 vccd1
+ _13650_/D sky130_fd_sc_hd__o221a_1
XFILLER_115_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _08792_/A vssd1 vssd1 vccd1 vccd1 _08767_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07718_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07718_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08698_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08698_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _14240_/Q _07644_/X _07428_/X _07646_/X _07640_/X vssd1 vssd1 vccd1 vccd1
+ _14240_/D sky130_fd_sc_hd__o221a_1
XPHY_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10660_ _13984_/Q vssd1 vssd1 vccd1 vccd1 _10660_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09319_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10591_ _13585_/Q vssd1 vssd1 vccd1 vccd1 _10591_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12330_ _13196_/Q _12329_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12330_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12261_ _12047_/Y _13362_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14000_ _14110_/CLK _14000_/D vssd1 vssd1 vccd1 vccd1 _14000_/Q sky130_fd_sc_hd__dfxtp_1
X_11212_ _14190_/Q vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12192_ vssd1 vssd1 vccd1 vccd1 _12192_/HI _12192_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11143_ _14384_/Q vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11074_ _11072_/Y _10987_/X _11073_/Y _10989_/X vssd1 vssd1 vccd1 vccd1 _11074_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput120 la_data_in[58] vssd1 vssd1 vccd1 vccd1 _06536_/A sky130_fd_sc_hd__buf_2
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput131 la_data_in[68] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__buf_1
XPHY_7152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10025_ _10025_/A vssd1 vssd1 vccd1 vccd1 _10026_/B sky130_fd_sc_hd__inv_2
Xinput142 la_data_in[78] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__buf_1
XFILLER_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput153 la_data_in[88] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_1
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 la_data_in[98] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_1
XPHY_7185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 la_oenb[107] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__buf_1
XFILLER_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput186 la_oenb[117] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_hd__buf_1
XPHY_6462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput197 la_oenb[127] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_1
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11976_ _14324_/Q vssd1 vssd1 vccd1 vccd1 _11976_/Y sky130_fd_sc_hd__inv_2
XPHY_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13715_ _14188_/CLK _13715_/D vssd1 vssd1 vccd1 vccd1 _13715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10927_ _11401_/A vssd1 vssd1 vccd1 vccd1 _10927_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13646_ _14139_/CLK _13646_/D vssd1 vssd1 vccd1 vccd1 _13646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10858_ _10848_/Y _10702_/X _10851_/X _10854_/X _10857_/X vssd1 vssd1 vccd1 vccd1
+ _10880_/C sky130_fd_sc_hd__o2111a_4
XFILLER_53_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13577_ _14130_/CLK _13577_/D vssd1 vssd1 vccd1 vccd1 _13577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10784_/Y _10735_/X _10785_/Y _10737_/X _10788_/X vssd1 vssd1 vccd1 vccd1
+ _10796_/C sky130_fd_sc_hd__o221a_1
XFILLER_160_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12528_ _13372_/Q _10035_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12528_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12459_ _12458_/X _06930_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12459_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput605 _13262_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _14130_/CLK _14129_/D vssd1 vssd1 vccd1 vccd1 _14129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06951_ _06954_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _14575_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09670_ _06897_/A _14581_/Q _14589_/Q _06927_/Y vssd1 vssd1 vccd1 vccd1 _09671_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_45_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06882_ _06976_/A vssd1 vssd1 vccd1 vccd1 _06958_/A sky130_fd_sc_hd__buf_2
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08621_ _13764_/Q _08618_/X _08527_/X _08619_/X _08620_/X vssd1 vssd1 vccd1 vccd1
+ _13764_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08552_ _08552_/A vssd1 vssd1 vccd1 vccd1 _08552_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07503_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07503_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08483_ _08745_/A _10207_/A vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__or2_2
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07365_ _08153_/A vssd1 vssd1 vccd1 vccd1 _07365_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_148_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09104_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07296_ _14409_/Q _07290_/X _06834_/X _07291_/X _07295_/X vssd1 vssd1 vccd1 vccd1
+ _14409_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09035_ _09035_/A vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__buf_4
XFILLER_178_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _09937_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09868_ _13300_/Q vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__inv_2
XFILLER_189_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08819_ _08877_/A vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_189_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09799_ _13344_/Q _09794_/Y _09801_/B vssd1 vssd1 vccd1 vccd1 _09799_/X sky130_fd_sc_hd__o21a_1
XPHY_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11830_/A vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11761_ _13571_/Q _11664_/X _13812_/Q _11665_/X vssd1 vssd1 vccd1 vccd1 _11761_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _14094_/CLK _13500_/D vssd1 vssd1 vccd1 vccd1 _13500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10708_/Y _10709_/X _10710_/Y _10711_/X vssd1 vssd1 vccd1 vccd1 _10712_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14481_/CLK _14480_/D vssd1 vssd1 vccd1 vccd1 _14480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11692_ _13491_/Q vssd1 vssd1 vccd1 vccd1 _11692_/Y sky130_fd_sc_hd__inv_2
XPHY_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13431_ _14143_/CLK _13431_/D vssd1 vssd1 vccd1 vccd1 _13431_/Q sky130_fd_sc_hd__dfxtp_1
X_10643_ _10624_/X _10643_/B _10643_/C _10643_/D vssd1 vssd1 vccd1 vccd1 _10644_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13362_ _14639_/CLK _13362_/D vssd1 vssd1 vccd1 vccd1 _13362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10574_ _10572_/Y _10448_/X _10573_/Y _10451_/X vssd1 vssd1 vccd1 vccd1 _10574_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12313_ _10685_/Y _14530_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12313_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13293_ _13877_/CLK _13293_/D vssd1 vssd1 vccd1 vccd1 _13293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12244_ _12244_/A vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12175_ vssd1 vssd1 vccd1 vccd1 _12175_/HI _12175_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ _14228_/Q _10933_/X _14423_/Q _10935_/X _11125_/X vssd1 vssd1 vccd1 vccd1
+ _11159_/B sky130_fd_sc_hd__a221oi_2
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11057_ _13208_/Q _11013_/X _14031_/Q _10957_/X _11056_/X vssd1 vssd1 vccd1 vccd1
+ _11057_/X sky130_fd_sc_hd__a221o_4
XFILLER_81_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10008_ _13375_/Q _10008_/B vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11959_ _13895_/Q vssd1 vssd1 vccd1 vccd1 _11959_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13629_ _14071_/CLK _13629_/D vssd1 vssd1 vccd1 vccd1 _13629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _14487_/Q _07144_/X _06834_/X _07145_/X _07147_/X vssd1 vssd1 vccd1 vccd1
+ _14487_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07081_ _14523_/Q _07014_/A _06845_/X _07017_/A _07079_/X vssd1 vssd1 vccd1 vccd1
+ _14523_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput402 _12202_/X vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__clkbuf_2
Xoutput413 _12092_/LO vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput424 _12240_/A vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput435 _12232_/A vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__clkbuf_2
Xoutput446 _12098_/LO vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput457 _12244_/X vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput468 _10129_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput479 _12112_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07983_ _08000_/A vssd1 vssd1 vccd1 vccd1 _07983_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ _09641_/Y _09721_/X _09641_/Y _09721_/X vssd1 vssd1 vccd1 vccd1 _09722_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06934_ _06919_/X _12303_/X _06933_/Y _06921_/X vssd1 vssd1 vccd1 vccd1 _06935_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09653_ _09644_/X _09652_/X _09644_/X _09652_/X vssd1 vssd1 vccd1 vccd1 _09653_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06865_ _06865_/A vssd1 vssd1 vccd1 vccd1 _06865_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08604_ _13774_/Q _08599_/X _08501_/X _08601_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _13774_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09584_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06796_ _08155_/A vssd1 vssd1 vccd1 vccd1 _06796_/X sky130_fd_sc_hd__buf_4
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ _13800_/Q _08526_/X _08534_/X _08528_/X _08524_/X vssd1 vssd1 vccd1 vccd1
+ _13800_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _13829_/Q _08460_/X _08169_/X _08461_/X _08465_/X vssd1 vssd1 vccd1 vccd1
+ _13829_/D sky130_fd_sc_hd__o221a_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _14363_/Q _07411_/X _07311_/X _07414_/X _07415_/X vssd1 vssd1 vccd1 vccd1
+ _14363_/D sky130_fd_sc_hd__o221a_1
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08397_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07279_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07279_/X sky130_fd_sc_hd__buf_2
X_09018_ _13565_/Q _09014_/X _08922_/X _09015_/X _09011_/X vssd1 vssd1 vccd1 vccd1
+ _13565_/D sky130_fd_sc_hd__o221a_1
XFILLER_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10290_ _10285_/Y _10228_/X _10286_/Y _10231_/X _10289_/X vssd1 vssd1 vccd1 vccd1
+ _10297_/C sky130_fd_sc_hd__o221a_1
XFILLER_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13980_ _14100_/CLK _13980_/D vssd1 vssd1 vccd1 vccd1 _13980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ _12545_/X _12930_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12931_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12862_ _12526_/X _12861_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XPHY_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14601_ _14637_/CLK _14601_/D vssd1 vssd1 vccd1 vccd1 _14601_/Q sky130_fd_sc_hd__dfxtp_1
X_11813_ _14281_/Q vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__inv_2
XPHY_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12793_ _09537_/X _12792_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12793_/X sky130_fd_sc_hd__mux2_1
XPHY_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14611_/CLK _14532_/D vssd1 vssd1 vccd1 vccd1 _14532_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11744_ _13649_/Q vssd1 vssd1 vccd1 vccd1 _11744_/Y sky130_fd_sc_hd__inv_2
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14595_/CLK _14463_/D vssd1 vssd1 vccd1 vccd1 _14463_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11675_/A vssd1 vssd1 vccd1 vccd1 _11675_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _14178_/CLK _13414_/D vssd1 vssd1 vccd1 vccd1 _13414_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10626_ _14334_/Q vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__inv_2
X_14394_ _14629_/CLK _14394_/D vssd1 vssd1 vccd1 vccd1 _14394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13345_ _14538_/CLK _13345_/D vssd1 vssd1 vccd1 vccd1 _13345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10557_ _14449_/Q vssd1 vssd1 vccd1 vccd1 _10557_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13276_ _13370_/CLK _13276_/D vssd1 vssd1 vccd1 vccd1 _13276_/Q sky130_fd_sc_hd__dfxtp_4
X_10488_ _10482_/Y _10484_/X _10485_/Y _10487_/X vssd1 vssd1 vccd1 vccd1 _10488_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12227_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ vssd1 vssd1 vccd1 vccd1 _12158_/HI _12158_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11109_ _11107_/Y _10977_/X _11108_/Y _10979_/X vssd1 vssd1 vccd1 vccd1 _11109_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12089_ vssd1 vssd1 vccd1 vccd1 _12089_/HI _12089_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06650_ _06643_/X _06649_/X _06643_/X _06649_/X vssd1 vssd1 vccd1 vccd1 _06829_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06581_ _06566_/X _06580_/Y _06566_/X _06580_/Y vssd1 vssd1 vccd1 vccd1 _06581_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08320_ _13910_/Q _08318_/X _08162_/X _08319_/X _08313_/X vssd1 vssd1 vccd1 vccd1
+ _13910_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08251_ _13948_/Q _08246_/X _08165_/X _08247_/X _08249_/X vssd1 vssd1 vccd1 vccd1
+ _13948_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07202_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08182_ _13980_/Q _08174_/X _08181_/X _08176_/X _08172_/X vssd1 vssd1 vccd1 vccd1
+ _13980_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07133_ _14498_/Q _07127_/X _06796_/X _07128_/X _07131_/X vssd1 vssd1 vccd1 vccd1
+ _14498_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07064_ _14534_/Q _07061_/X _06807_/X _07062_/X _07063_/X vssd1 vssd1 vccd1 vccd1
+ _14534_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07966_ _08008_/A vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__buf_6
XFILLER_102_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09705_ _09684_/A _09704_/X _09684_/A _09704_/X vssd1 vssd1 vccd1 vccd1 _09705_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_210_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06917_ _06917_/A _06917_/B vssd1 vssd1 vccd1 vccd1 _14584_/D sky130_fd_sc_hd__nor2_1
X_07897_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07897_/X sky130_fd_sc_hd__buf_2
XFILLER_99_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _06957_/Y _14569_/Q _14573_/Q _06970_/Y vssd1 vssd1 vccd1 vccd1 _09637_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06848_ _14600_/Q _06530_/A _06716_/X _08190_/A _06838_/X vssd1 vssd1 vccd1 vccd1
+ _14600_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09567_ _09573_/A _12358_/X vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__and2_1
XFILLER_58_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06779_ _14620_/Q _06769_/X _06778_/X _06772_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _14620_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08518_ _13807_/Q _08513_/X _08517_/X _08515_/X _08511_/X vssd1 vssd1 vccd1 vccd1
+ _13807_/D sky130_fd_sc_hd__o221a_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _13263_/Q _09493_/X _12258_/X _09494_/X vssd1 vssd1 vccd1 vccd1 _13263_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08449_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11460_ _14468_/Q vssd1 vssd1 vccd1 vccd1 _11460_/Y sky130_fd_sc_hd__inv_2
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10411_ _14174_/Q vssd1 vssd1 vccd1 vccd1 _10411_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _14467_/Q vssd1 vssd1 vccd1 vccd1 _11391_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13130_ _13129_/X _12643_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ _13425_/Q vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13061_ _12610_/X _13060_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10273_ _10271_/Y _10195_/X _10272_/Y _10198_/X vssd1 vssd1 vccd1 vccd1 _10273_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12012_ _14364_/Q vssd1 vssd1 vccd1 vccd1 _12012_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13963_ _14110_/CLK _13963_/D vssd1 vssd1 vccd1 vccd1 _13963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12914_ _12539_/X _12913_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12914_/X sky130_fd_sc_hd__mux2_1
X_13894_ _14130_/CLK _13894_/D vssd1 vssd1 vccd1 vccd1 _13894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12845_ _12522_/X _12844_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12776_ _09524_/X input350/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__mux2_1
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _14318_/Q vssd1 vssd1 vccd1 vccd1 _11727_/Y sky130_fd_sc_hd__inv_2
X_14515_ _14633_/CLK _14515_/D vssd1 vssd1 vccd1 vccd1 _14515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11658_/A vssd1 vssd1 vccd1 vccd1 _11658_/X sky130_fd_sc_hd__clkbuf_2
X_14446_ _14481_/CLK _14446_/D vssd1 vssd1 vccd1 vccd1 _14446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _10604_/Y _10425_/X _10605_/Y _10428_/X _10608_/X vssd1 vssd1 vccd1 vccd1
+ _10644_/A sky130_fd_sc_hd__o221a_2
XFILLER_102_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _14627_/CLK _14377_/D vssd1 vssd1 vccd1 vccd1 _14377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11589_ _11570_/X _11589_/B _11589_/C _11589_/D vssd1 vssd1 vccd1 vccd1 _11590_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_89_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13328_ _13877_/CLK _13328_/D vssd1 vssd1 vccd1 vccd1 _13328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13259_ _14639_/CLK _13259_/D vssd1 vssd1 vccd1 vccd1 _13259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07856_/A sky130_fd_sc_hd__buf_6
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater702 _13109_/S vssd1 vssd1 vccd1 vccd1 _13085_/S sky130_fd_sc_hd__buf_4
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07751_ _08142_/A vssd1 vssd1 vccd1 vccd1 _07751_/X sky130_fd_sc_hd__buf_6
XFILLER_113_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06702_ _06701_/X _06667_/Y _06701_/X _06667_/Y vssd1 vssd1 vccd1 vccd1 _09035_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07682_ _14221_/Q _07679_/X _07377_/X _07680_/X _07676_/X vssd1 vssd1 vccd1 vccd1
+ _14221_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09421_ _09445_/A vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06633_ _06593_/Y _08925_/A _08914_/A _06564_/Y vssd1 vssd1 vccd1 vccd1 _06633_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09352_ _09352_/A vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06564_ _06565_/A vssd1 vssd1 vccd1 vccd1 _06564_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08303_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09283_ _13417_/Q _09275_/X _07714_/A _09277_/X _09280_/X vssd1 vssd1 vccd1 vccd1
+ _13417_/D sky130_fd_sc_hd__o221a_1
X_06495_ _06495_/A _06495_/B _06495_/C _06495_/D vssd1 vssd1 vccd1 vccd1 _06498_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_181_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _13957_/Q _08229_/X _08142_/X _08230_/X _08231_/X vssd1 vssd1 vccd1 vccd1
+ _13957_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08165_ _08165_/A vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__buf_4
XFILLER_14_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07116_ _14508_/Q _07111_/X _06760_/X _07112_/X _07114_/X vssd1 vssd1 vccd1 vccd1
+ _14508_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08096_ _08176_/A vssd1 vssd1 vccd1 vccd1 _08097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07047_ _14544_/Q _07044_/X _06771_/X _07045_/X _07046_/X vssd1 vssd1 vccd1 vccd1
+ _14544_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _13575_/Q _08993_/X _08825_/X _08995_/X _08986_/X vssd1 vssd1 vccd1 vccd1
+ _13575_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ _14092_/Q _07882_/A _07876_/X _07884_/A _07946_/X vssd1 vssd1 vccd1 vccd1
+ _14092_/D sky130_fd_sc_hd__o221a_1
XPHY_6858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10960_ _13554_/Q _10958_/X _13795_/Q _10959_/X vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _09610_/Y _09618_/X _09610_/Y _09618_/X vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10891_ _13872_/Q vssd1 vssd1 vccd1 vccd1 _10891_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _09838_/Y _13329_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12561_ _09951_/X _13300_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__mux2_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11512_ _11510_/Y _11401_/X _11511_/Y _11403_/X vssd1 vssd1 vccd1 vccd1 _11512_/X
+ sky130_fd_sc_hd__o22a_2
X_14300_ _14305_/CLK _14300_/D vssd1 vssd1 vccd1 vccd1 _14300_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12492_ _12491_/X _06975_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__mux2_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14231_ _14595_/CLK _14231_/D vssd1 vssd1 vccd1 vccd1 _14231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11443_ _11434_/Y _11435_/X _11436_/Y _11437_/X _11442_/X vssd1 vssd1 vccd1 vccd1
+ _11464_/B sky130_fd_sc_hd__o221a_2
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14291_/CLK _14162_/D vssd1 vssd1 vccd1 vccd1 _14162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11374_ _13563_/Q _11194_/X _13804_/Q _11195_/X vssd1 vssd1 vccd1 vccd1 _11374_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13113_ _12635_/X _13112_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__mux2_1
X_10325_ _10323_/Y _10220_/X _10324_/Y _10223_/X vssd1 vssd1 vccd1 vccd1 _10325_/X
+ sky130_fd_sc_hd__o22a_1
X_14093_ _14094_/CLK _14093_/D vssd1 vssd1 vccd1 vccd1 _14093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13044_ _12602_/X input347/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13044_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10256_ _14054_/Q vssd1 vssd1 vccd1 vccd1 _10256_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10187_ _11653_/A vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__buf_2
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _14107_/CLK _13946_/D vssd1 vssd1 vccd1 vccd1 _13946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13877_ _13877_/CLK _13877_/D vssd1 vssd1 vccd1 vccd1 _13877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12828_ _12518_/X input336/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12759_ _09554_/X _12758_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13208_/D sky130_fd_sc_hd__mux2_1
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14429_ _14611_/CLK _14429_/D vssd1 vssd1 vccd1 vccd1 _14429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09970_ _13356_/Q _09970_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__nand2_1
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08921_ _13605_/Q _08916_/X _08920_/X _08918_/X _08910_/X vssd1 vssd1 vccd1 vccd1
+ _13605_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ _08868_/A vssd1 vssd1 vccd1 vccd1 _08852_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07803_ _07803_/A vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08783_ _08792_/A vssd1 vssd1 vccd1 vccd1 _08783_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07734_ _07772_/A vssd1 vssd1 vccd1 vccd1 _07734_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07665_ _14230_/Q _07661_/X _07354_/X _07662_/X _07658_/X vssd1 vssd1 vccd1 vccd1
+ _14230_/D sky130_fd_sc_hd__o221a_1
XFILLER_96_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09404_ _09407_/A _13099_/X vssd1 vssd1 vccd1 vccd1 _13331_/D sky130_fd_sc_hd__and2_1
XFILLER_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06616_ _06541_/Y _06553_/Y _06541_/A _06553_/A vssd1 vssd1 vccd1 vccd1 _06616_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07596_ _14267_/Q _07589_/X _07358_/X _07590_/X _07593_/X vssd1 vssd1 vccd1 vccd1
+ _14267_/D sky130_fd_sc_hd__o221a_1
XFILLER_209_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _13385_/Q _09275_/A _08188_/A _09277_/A _09330_/X vssd1 vssd1 vccd1 vccd1
+ _13385_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06547_ _08827_/A _06544_/Y _06545_/Y _08829_/A vssd1 vssd1 vccd1 vccd1 _06547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09266_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_178_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08217_ _08217_/A vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09197_ _13464_/Q _09135_/A _08981_/X _09137_/A _09196_/X vssd1 vssd1 vccd1 vccd1
+ _13464_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08148_ _13994_/Q _08136_/X _08146_/X _08138_/X _08147_/X vssd1 vssd1 vccd1 vccd1
+ _13994_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ _08079_/A vssd1 vssd1 vccd1 vccd1 _08079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10110_ _10145_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _12464_/S sky130_fd_sc_hd__or2_1
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _13837_/Q vssd1 vssd1 vccd1 vccd1 _11090_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _13362_/Q _09982_/B _09983_/A vssd1 vssd1 vccd1 vccd1 _10041_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput302 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _06502_/D sky130_fd_sc_hd__clkbuf_1
XPHY_7323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput313 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _06494_/B sky130_fd_sc_hd__clkbuf_1
XPHY_7334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput324 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _06507_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput335 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 input335/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput346 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 input346/X sky130_fd_sc_hd__clkbuf_8
XPHY_7367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput357 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input357/X sky130_fd_sc_hd__clkbuf_4
XPHY_7378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13800_ _14114_/CLK _13800_/D vssd1 vssd1 vccd1 vccd1 _13800_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ _13694_/Q vssd1 vssd1 vccd1 vccd1 _11992_/Y sky130_fd_sc_hd__inv_2
XPHY_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13731_ _14056_/CLK _13731_/D vssd1 vssd1 vccd1 vccd1 _13731_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _13873_/Q vssd1 vssd1 vccd1 vccd1 _10943_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13662_ _14047_/CLK _13662_/D vssd1 vssd1 vccd1 vccd1 _13662_/Q sky130_fd_sc_hd__dfxtp_1
X_10874_ _14144_/Q vssd1 vssd1 vccd1 vccd1 _10874_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ _09851_/Y _13322_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__mux2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _14188_/CLK _13593_/D vssd1 vssd1 vccd1 vccd1 _13593_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12544_ _09963_/X _13293_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _12474_/X _06952_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12475_/X sky130_fd_sc_hd__mux2_2
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14214_ _14291_/CLK _14214_/D vssd1 vssd1 vccd1 vccd1 _14214_/Q sky130_fd_sc_hd__dfxtp_1
X_11426_ _11426_/A vssd1 vssd1 vccd1 vccd1 _11426_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_6 _11035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _14146_/CLK _14145_/D vssd1 vssd1 vccd1 vccd1 _14145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11357_ _13680_/Q vssd1 vssd1 vccd1 vccd1 _11357_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _13938_/Q vssd1 vssd1 vccd1 vccd1 _10308_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14076_ _14188_/CLK _14076_/D vssd1 vssd1 vccd1 vccd1 _14076_/Q sky130_fd_sc_hd__dfxtp_1
X_11288_ _13997_/Q vssd1 vssd1 vccd1 vccd1 _11288_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13027_ _12592_/X _13026_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__mux2_1
X_10239_ _10226_/Y _10228_/X _10229_/Y _10231_/X _10238_/X vssd1 vssd1 vccd1 vccd1
+ _10254_/C sky130_fd_sc_hd__o221a_1
XFILLER_140_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _14139_/CLK _13929_/D vssd1 vssd1 vccd1 vccd1 _13929_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07450_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07381_ _08169_/A vssd1 vssd1 vccd1 vccd1 _07381_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09120_ _09120_/A vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _09051_/A vssd1 vssd1 vccd1 vccd1 _09051_/X sky130_fd_sc_hd__buf_4
XFILLER_175_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08002_ _14065_/Q _07999_/X _07774_/X _08000_/X _07995_/X vssd1 vssd1 vccd1 vccd1
+ _14065_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09953_ _09895_/A _09895_/B _09952_/Y vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08956_/A sky130_fd_sc_hd__buf_4
XFILLER_98_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09884_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__or2_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08835_ _08869_/A vssd1 vssd1 vccd1 vccd1 _08835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _13685_/Q _08758_/X _08510_/X _08760_/X _08761_/X vssd1 vssd1 vccd1 vccd1
+ _13685_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07717_ _07783_/A vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__buf_4
XPHY_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08697_ _13724_/Q _08687_/X _08510_/X _08689_/X _08696_/X vssd1 vssd1 vccd1 vccd1
+ _13724_/D sky130_fd_sc_hd__o221a_1
XPHY_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ _14241_/Q _07644_/X _07327_/X _07646_/X _07640_/X vssd1 vssd1 vccd1 vccd1
+ _14241_/D sky130_fd_sc_hd__o221a_1
XPHY_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07579_ _14277_/Q _07571_/X _07332_/X _07573_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _14277_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09318_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09318_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ _14294_/Q vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09249_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12260_ _12046_/Y _13361_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ _11447_/A vssd1 vssd1 vccd1 vccd1 _11211_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12191_ vssd1 vssd1 vccd1 vccd1 _12191_/HI _12191_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11142_ _14618_/Q vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11073_ _14460_/Q vssd1 vssd1 vccd1 vccd1 _11073_/Y sky130_fd_sc_hd__inv_2
XPHY_7120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 la_data_in[49] vssd1 vssd1 vccd1 vccd1 _06609_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput121 la_data_in[59] vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__buf_2
XFILLER_209_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10024_ _13380_/Q _10023_/B _10025_/A vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__o21a_1
Xinput132 la_data_in[69] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__buf_1
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput143 la_data_in[79] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__buf_1
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput154 la_data_in[89] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__buf_1
XFILLER_23_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput165 la_data_in[99] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_1
XPHY_7186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 la_oenb[108] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_hd__buf_1
XPHY_7197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput187 la_oenb[118] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_hd__buf_1
XPHY_6463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput198 la_oenb[12] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__buf_1
XFILLER_40_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _11970_/Y _10214_/A _11971_/Y _10217_/A _11974_/X vssd1 vssd1 vccd1 vccd1
+ _11988_/B sky130_fd_sc_hd__o221a_4
XPHY_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13714_ _14188_/CLK _13714_/D vssd1 vssd1 vccd1 vccd1 _13714_/Q sky130_fd_sc_hd__dfxtp_1
X_10926_ _13671_/Q vssd1 vssd1 vccd1 vccd1 _10926_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13645_ _14143_/CLK _13645_/D vssd1 vssd1 vccd1 vccd1 _13645_/Q sky130_fd_sc_hd__dfxtp_1
X_10857_ _10855_/Y _10714_/X _10856_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _10857_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _14130_/CLK _13576_/D vssd1 vssd1 vccd1 vccd1 _13576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10788_ _10786_/Y _10739_/X _10787_/Y _10741_/X vssd1 vssd1 vccd1 vccd1 _10788_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12527_ _13373_/Q _10036_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12458_ _12509_/X _06930_/Y _12458_/S vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput606 _13263_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _13408_/Q _11278_/X _13720_/Q _11408_/X vssd1 vssd1 vccd1 vccd1 _11409_/X
+ sky130_fd_sc_hd__a22o_2
X_12389_ _13208_/Q _06602_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _14130_/CLK _14128_/D vssd1 vssd1 vccd1 vccd1 _14128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06950_ _06937_/X _12307_/X _06949_/Y _06939_/X vssd1 vssd1 vccd1 vccd1 _06951_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14059_ _14139_/CLK _14059_/D vssd1 vssd1 vccd1 vccd1 _14059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06881_ _14593_/Q vssd1 vssd1 vccd1 vccd1 _06881_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08620_ _08637_/A vssd1 vssd1 vccd1 vccd1 _08620_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _13794_/Q _08540_/X _08549_/X _08542_/X _08550_/X vssd1 vssd1 vccd1 vccd1
+ _13794_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07502_ _14320_/Q _07499_/X _07323_/X _07501_/X _07493_/X vssd1 vssd1 vccd1 vccd1
+ _14320_/D sky130_fd_sc_hd__o221a_1
X_08482_ _08989_/A _08482_/B _08989_/C _08482_/D vssd1 vssd1 vccd1 vccd1 _10207_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_1_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07433_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07433_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07364_ _14383_/Q _07361_/X _07362_/X _07363_/X _07359_/X vssd1 vssd1 vccd1 vccd1
+ _14383_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09103_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09103_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07295_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09034_ _13555_/Q _09030_/X _08950_/X _09031_/X _09027_/X vssd1 vssd1 vccd1 vccd1
+ _13555_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09936_ _13306_/Q _09934_/Y _09901_/B vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09867_ _13301_/Q vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__inv_2
XFILLER_150_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08818_ _08818_/A vssd1 vssd1 vccd1 vccd1 _08818_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__or2_1
XFILLER_189_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _13272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _08801_/A vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__clkbuf_2
XPHY_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11760_ _11750_/Y _11646_/X _11753_/X _11756_/X _11759_/X vssd1 vssd1 vccd1 vccd1
+ _11782_/C sky130_fd_sc_hd__o2111a_4
XPHY_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _11421_/A vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _11691_/A vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__buf_2
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _10637_/Y _10506_/X _10638_/Y _10509_/X _10641_/X vssd1 vssd1 vccd1 vccd1
+ _10643_/D sky130_fd_sc_hd__o221a_1
X_13430_ _14139_/CLK _13430_/D vssd1 vssd1 vccd1 vccd1 _13430_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13361_ _14639_/CLK _13361_/D vssd1 vssd1 vccd1 vccd1 _13361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10573_ _13865_/Q vssd1 vssd1 vccd1 vccd1 _10573_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12312_ _10755_/Y _14531_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12312_/X sky130_fd_sc_hd__mux2_2
XFILLER_196_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13292_ _13877_/CLK _13292_/D vssd1 vssd1 vccd1 vccd1 _13292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12243_ _12243_/A vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12174_ vssd1 vssd1 vccd1 vccd1 _12174_/HI _12174_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11125_ _13402_/Q _11042_/X _13714_/Q _10936_/X vssd1 vssd1 vccd1 vccd1 _11125_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11056_ _13556_/Q _10958_/X _13797_/Q _10959_/X vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _10008_/B sky130_fd_sc_hd__inv_2
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _13778_/Q vssd1 vssd1 vccd1 vccd1 _11958_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10909_ _13592_/Q vssd1 vssd1 vccd1 vccd1 _10909_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11889_ _14361_/Q vssd1 vssd1 vccd1 vccd1 _11889_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13628_ _14071_/CLK _13628_/D vssd1 vssd1 vccd1 vccd1 _13628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13559_ _14114_/CLK _13559_/D vssd1 vssd1 vccd1 vccd1 _13559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07080_ _14524_/Q _07014_/A _06843_/B _07017_/A _07079_/X vssd1 vssd1 vccd1 vccd1
+ _14524_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput403 _12203_/X vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput414 _12093_/LO vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput425 _12241_/A vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput436 _12233_/A vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput447 _12099_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput458 _12109_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput469 _12110_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07982_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07982_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06933_ _14579_/Q vssd1 vssd1 vccd1 vccd1 _06933_/Y sky130_fd_sc_hd__inv_2
X_09721_ _14576_/Q _14575_/Q _06946_/Y _06949_/Y vssd1 vssd1 vccd1 vccd1 _09721_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09652_ _06989_/X _09651_/X _06989_/X _09651_/X vssd1 vssd1 vccd1 vccd1 _09652_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06864_ _14597_/Q vssd1 vssd1 vccd1 vccd1 _06865_/A sky130_fd_sc_hd__inv_2
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08603_ _08637_/A vssd1 vssd1 vccd1 vccd1 _08603_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09583_ _09583_/A vssd1 vssd1 vccd1 vccd1 _09583_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06795_ _08950_/A vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__buf_2
XFILLER_58_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _08940_/A vssd1 vssd1 vccd1 vccd1 _08534_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08465_/X sky130_fd_sc_hd__clkbuf_2
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ _14364_/Q _07411_/X _07412_/X _07414_/X _07415_/X vssd1 vssd1 vccd1 vccd1
+ _14364_/D sky130_fd_sc_hd__o221a_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08396_ _08396_/A vssd1 vssd1 vccd1 vccd1 _08396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07347_ _14389_/Q _07335_/X _07345_/X _07337_/X _07346_/X vssd1 vssd1 vccd1 vccd1
+ _14389_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07278_ _14420_/Q _07274_/X _06796_/X _07275_/X _07271_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/D sky130_fd_sc_hd__o221a_1
X_09017_ _13566_/Q _09014_/X _08920_/X _09015_/X _09011_/X vssd1 vssd1 vccd1 vccd1
+ _13566_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or2_1
XFILLER_154_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12930_ _12929_/X _12545_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12526_/X _12860_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14600_ _14637_/CLK _14600_/D vssd1 vssd1 vccd1 vccd1 _14600_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11812_ _14203_/Q vssd1 vssd1 vccd1 vccd1 _11812_/Y sky130_fd_sc_hd__inv_2
XPHY_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _09537_/X input346/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__mux2_1
XPHY_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14611_/CLK _14531_/D vssd1 vssd1 vccd1 vccd1 _14531_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13688_/Q vssd1 vssd1 vccd1 vccd1 _11743_/Y sky130_fd_sc_hd__inv_2
XPHY_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14462_ _14495_/CLK _14462_/D vssd1 vssd1 vccd1 vccd1 _14462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11674_ _14395_/Q vssd1 vssd1 vccd1 vccd1 _11674_/Y sky130_fd_sc_hd__inv_2
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _14178_/CLK _13413_/D vssd1 vssd1 vccd1 vccd1 _13413_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _14490_/Q vssd1 vssd1 vccd1 vccd1 _10625_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14393_ _14629_/CLK _14393_/D vssd1 vssd1 vccd1 vccd1 _14393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10556_ _13467_/Q vssd1 vssd1 vccd1 vccd1 _10556_/Y sky130_fd_sc_hd__inv_2
X_13344_ _14538_/CLK _13344_/D vssd1 vssd1 vccd1 vccd1 _13344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ _11441_/A vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__clkbuf_2
X_13275_ _13371_/CLK _13275_/D vssd1 vssd1 vccd1 vccd1 _13275_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_120_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12226_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ vssd1 vssd1 vccd1 vccd1 _12157_/HI _12157_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _14266_/Q vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12088_ vssd1 vssd1 vccd1 vccd1 _12088_/HI _12088_/LO sky130_fd_sc_hd__conb_1
XFILLER_209_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ _13634_/Q vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06580_ _06571_/X _06579_/X _06571_/X _06579_/X vssd1 vssd1 vccd1 vccd1 _06580_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08250_ _13949_/Q _08246_/X _08162_/X _08247_/X _08249_/X vssd1 vssd1 vccd1 vccd1
+ _13949_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07201_ _07209_/A vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08181_ _08181_/A vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__buf_4
XFILLER_146_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07132_ _14499_/Q _07127_/X _06793_/X _07128_/X _07131_/X vssd1 vssd1 vccd1 vccd1
+ _14499_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07063_ _07071_/A vssd1 vssd1 vccd1 vccd1 _07063_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07965_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07965_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09704_ _09699_/X _09703_/X _09699_/X _09703_/X vssd1 vssd1 vccd1 vccd1 _09704_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06916_ _06901_/X _12298_/X _06915_/Y _06903_/X vssd1 vssd1 vccd1 vccd1 _06917_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07896_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09635_ _09631_/X _09634_/X _09631_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _09635_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06847_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08190_/A sky130_fd_sc_hd__buf_4
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09566_ _09557_/X _09565_/X _13268_/Q _09558_/X vssd1 vssd1 vccd1 vccd1 _13236_/D
+ sky130_fd_sc_hd__o22a_1
X_06778_ _08142_/A vssd1 vssd1 vccd1 vccd1 _06778_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08517_ _08920_/A vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _13264_/Q _09493_/X _12259_/X _09494_/X vssd1 vssd1 vccd1 vccd1 _13264_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08448_ _13840_/Q _08444_/X _08142_/X _08445_/X _08441_/X vssd1 vssd1 vccd1 vccd1
+ _13840_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08379_ _08388_/A vssd1 vssd1 vccd1 vccd1 _08379_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10410_ _13582_/Q vssd1 vssd1 vccd1 vccd1 _10410_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _13485_/Q vssd1 vssd1 vccd1 vccd1 _11390_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10341_ _14056_/Q vssd1 vssd1 vccd1 vccd1 _10341_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ _12610_/X input357/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__mux2_1
X_10272_ _13501_/Q vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _14520_/Q vssd1 vssd1 vccd1 vccd1 _12011_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13962_ _14110_/CLK _13962_/D vssd1 vssd1 vccd1 vccd1 _13962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12913_ _12539_/X _12912_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__mux2_1
X_13893_ _14130_/CLK _13893_/D vssd1 vssd1 vccd1 vccd1 _13893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12844_ _12522_/X input332/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12775_ _09522_/X _12774_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13220_/D sky130_fd_sc_hd__mux2_1
XFILLER_37_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14633_/CLK _14514_/D vssd1 vssd1 vccd1 vccd1 _14514_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11721_/Y _11669_/X _11722_/Y _11671_/X _11725_/X vssd1 vssd1 vccd1 vccd1
+ _11739_/B sky130_fd_sc_hd__o221a_2
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14445_ _14481_/CLK _14445_/D vssd1 vssd1 vccd1 vccd1 _14445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _14005_/Q vssd1 vssd1 vccd1 vccd1 _11657_/Y sky130_fd_sc_hd__inv_2
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ _10606_/Y _10431_/X _10607_/Y _10434_/X vssd1 vssd1 vccd1 vccd1 _10608_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14627_/CLK _14376_/D vssd1 vssd1 vccd1 vccd1 _14376_/Q sky130_fd_sc_hd__dfxtp_1
X_11588_ _11583_/Y _11455_/X _11584_/Y _11457_/X _11587_/X vssd1 vssd1 vccd1 vccd1
+ _11589_/D sky130_fd_sc_hd__o221a_1
XFILLER_102_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13327_ _13877_/CLK _13327_/D vssd1 vssd1 vccd1 vccd1 _13327_/Q sky130_fd_sc_hd__dfxtp_1
X_10539_ _11013_/A vssd1 vssd1 vccd1 vccd1 _10539_/X sky130_fd_sc_hd__buf_2
XFILLER_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13258_ _14639_/CLK _13258_/D vssd1 vssd1 vccd1 vccd1 _13258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _06865_/X _06858_/Y _06872_/Y _06869_/X _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13189_/X sky130_fd_sc_hd__mux4_2
XFILLER_83_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater703 _13113_/S vssd1 vssd1 vccd1 vccd1 _13109_/S sky130_fd_sc_hd__buf_8
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07750_ _14192_/Q _07745_/X _07749_/X _07747_/X _07743_/X vssd1 vssd1 vccd1 vccd1
+ _14192_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06701_ _06698_/X _06700_/X _06698_/X _06700_/X vssd1 vssd1 vccd1 vccd1 _06701_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07681_ _14222_/Q _07679_/X _07374_/X _07680_/X _07676_/X vssd1 vssd1 vccd1 vccd1
+ _14222_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09420_ _09509_/A vssd1 vssd1 vccd1 vccd1 _09445_/A sky130_fd_sc_hd__buf_4
X_06632_ _06632_/A vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09351_ _09351_/A _12867_/X vssd1 vssd1 vccd1 vccd1 _13373_/D sky130_fd_sc_hd__and2_1
X_06563_ _06562_/A _06561_/Y _06562_/Y _06561_/A vssd1 vssd1 vccd1 vccd1 _06563_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08302_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08302_/X sky130_fd_sc_hd__clkbuf_2
X_09282_ _13418_/Q _09275_/X _07712_/A _09277_/X _09280_/X vssd1 vssd1 vccd1 vccd1
+ _13418_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06494_ _06494_/A _06494_/B _06494_/C _06494_/D vssd1 vssd1 vccd1 vccd1 _06498_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08233_ _13958_/Q _08229_/X _08140_/X _08230_/X _08231_/X vssd1 vssd1 vccd1 vccd1
+ _13958_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08164_ _13988_/Q _08161_/X _08162_/X _08163_/X _08159_/X vssd1 vssd1 vccd1 vccd1
+ _13988_/D sky130_fd_sc_hd__o221a_1
XFILLER_181_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07115_ _14509_/Q _07111_/X _06757_/X _07112_/X _07114_/X vssd1 vssd1 vccd1 vccd1
+ _14509_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _08095_/A vssd1 vssd1 vccd1 vccd1 _08095_/X sky130_fd_sc_hd__buf_2
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07046_ _07071_/A vssd1 vssd1 vccd1 vccd1 _07046_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ _13576_/Q _08993_/X _08822_/X _08995_/X _08986_/X vssd1 vssd1 vccd1 vccd1
+ _13576_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _14093_/Q _07882_/A _07800_/X _07884_/A _07946_/X vssd1 vssd1 vccd1 vccd1
+ _14093_/D sky130_fd_sc_hd__o221a_1
XPHY_6848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07879_ _07952_/A _11655_/A vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__or2_2
XFILLER_186_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09618_ _09616_/X _09617_/X _09616_/X _09617_/X vssd1 vssd1 vccd1 vccd1 _09618_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _13755_/Q vssd1 vssd1 vccd1 vccd1 _10890_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ _09588_/A vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__buf_1
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ _13301_/Q _12559_/X input39/X vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__mux2_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11511_ _13644_/Q vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12491_ _12509_/X _06975_/Y _12491_/S vssd1 vssd1 vccd1 vccd1 _12491_/X sky130_fd_sc_hd__mux2_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _14595_/CLK _14230_/D vssd1 vssd1 vccd1 vccd1 _14230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11442_ _11438_/Y _11439_/X _11440_/Y _11441_/X vssd1 vssd1 vccd1 vccd1 _11442_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14161_ _14291_/CLK _14161_/D vssd1 vssd1 vccd1 vccd1 _14161_/Q sky130_fd_sc_hd__dfxtp_1
X_11373_ _11363_/Y _11176_/X _11366_/X _11369_/X _11372_/X vssd1 vssd1 vccd1 vccd1
+ _11395_/C sky130_fd_sc_hd__o2111a_4
XFILLER_193_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10324_ _14367_/Q vssd1 vssd1 vccd1 vccd1 _10324_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13112_ _12635_/X input360/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14095_/CLK _14092_/D vssd1 vssd1 vccd1 vccd1 _14092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10255_ _10255_/A _10255_/B _10255_/C _10255_/D vssd1 vssd1 vccd1 vccd1 _10255_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_4_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _12600_/X _13042_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10186_ _13819_/Q vssd1 vssd1 vccd1 vccd1 _10186_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13945_ _14107_/CLK _13945_/D vssd1 vssd1 vccd1 vccd1 _13945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _13877_/CLK _13876_/D vssd1 vssd1 vccd1 vccd1 _13876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12827_ _10048_/X _12826_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12758_ _09554_/X _12757_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__mux2_1
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11709_ _13772_/Q vssd1 vssd1 vccd1 vccd1 _11709_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _09593_/X _12688_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12689_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _14611_/CLK _14428_/D vssd1 vssd1 vccd1 vccd1 _14428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14359_ _14629_/CLK _14359_/D vssd1 vssd1 vccd1 vccd1 _14359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _08920_/A vssd1 vssd1 vccd1 vccd1 _08920_/X sky130_fd_sc_hd__buf_6
XFILLER_83_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08851_ _13641_/Q _08844_/X _08523_/X _08845_/X _08847_/X vssd1 vssd1 vccd1 vccd1
+ _13641_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07802_ _14170_/Q _07704_/A _07480_/X _07706_/A _07794_/X vssd1 vssd1 vccd1 vccd1
+ _14170_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08782_ _13675_/Q _08775_/X _08536_/X _08776_/X _08777_/X vssd1 vssd1 vccd1 vccd1
+ _13675_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07733_ _08123_/A vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__buf_4
XFILLER_96_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07664_ _14231_/Q _07661_/X _07352_/X _07662_/X _07658_/X vssd1 vssd1 vccd1 vccd1
+ _14231_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09407_/A _13095_/X vssd1 vssd1 vccd1 vccd1 _13332_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06615_ _08942_/A _06603_/A _06614_/Y _06603_/Y vssd1 vssd1 vccd1 vccd1 _06615_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07595_ _14268_/Q _07589_/X _07356_/X _07590_/X _07593_/X vssd1 vssd1 vccd1 vccd1
+ _14268_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09334_ _13386_/Q _09275_/A _08186_/A _09277_/A _09330_/X vssd1 vssd1 vccd1 vccd1
+ _13386_/D sky130_fd_sc_hd__o221a_1
X_06546_ _06546_/A vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__buf_4
XFILLER_209_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09265_ _13425_/Q _09205_/A _08981_/X _09207_/A _09260_/X vssd1 vssd1 vccd1 vccd1
+ _13425_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _13968_/Q _08211_/X _08114_/X _08213_/X _08214_/X vssd1 vssd1 vccd1 vccd1
+ _13968_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09196_ _09219_/A vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__buf_2
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _08184_/A vssd1 vssd1 vccd1 vccd1 _08147_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08078_ _08078_/A vssd1 vssd1 vccd1 vccd1 _08078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07029_ _14554_/Q _07025_/X _06735_/X _07027_/X _07028_/X vssd1 vssd1 vccd1 vccd1
+ _14554_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _13361_/Q _09980_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _10040_/X sky130_fd_sc_hd__o21a_1
XPHY_7313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput303 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _06502_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput314 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _06494_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput325 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _06507_/C sky130_fd_sc_hd__clkbuf_1
XPHY_7346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput336 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 input336/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput347 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 input347/X sky130_fd_sc_hd__clkbuf_8
XPHY_7368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput358 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input358/X sky130_fd_sc_hd__clkbuf_4
XPHY_7379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ _13460_/Q vssd1 vssd1 vccd1 vccd1 _11991_/Y sky130_fd_sc_hd__inv_2
XPHY_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _14056_/CLK _13730_/D vssd1 vssd1 vccd1 vccd1 _13730_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10942_ _11414_/A vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13661_ _14047_/CLK _13661_/D vssd1 vssd1 vccd1 vccd1 _13661_/Q sky130_fd_sc_hd__dfxtp_1
X_10873_ _13910_/Q vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _13323_/Q _12611_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12612_/X sky130_fd_sc_hd__mux2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _14188_/CLK _13592_/D vssd1 vssd1 vccd1 vccd1 _13592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12543_ _13294_/Q _12542_/X input39/X vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _12473_/X _06952_/Y _12486_/S vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _14291_/CLK _14213_/D vssd1 vssd1 vccd1 vccd1 _14213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11425_ _13525_/Q vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_7 _11077_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14144_ _14183_/CLK _14144_/D vssd1 vssd1 vccd1 vccd1 _14144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11356_ _13446_/Q vssd1 vssd1 vccd1 vccd1 _11356_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10307_ _14211_/Q _10164_/X _14406_/Q _10167_/X _10306_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/B sky130_fd_sc_hd__a221oi_2
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14075_ _14459_/CLK _14075_/D vssd1 vssd1 vccd1 vccd1 _14075_/Q sky130_fd_sc_hd__dfxtp_1
X_11287_ _11285_/Y _11183_/X _11286_/Y _11185_/X vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13026_ _13025_/X _12592_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10238_ _10232_/Y _10234_/X _10235_/Y _10237_/X vssd1 vssd1 vccd1 vccd1 _10238_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10169_ _11514_/A vssd1 vssd1 vccd1 vccd1 _11042_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _14139_/CLK _13928_/D vssd1 vssd1 vccd1 vccd1 _13928_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13859_ _14095_/CLK _13859_/D vssd1 vssd1 vccd1 vccd1 _13859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07380_ _14376_/Q _07373_/X _07379_/X _07375_/X _07371_/X vssd1 vssd1 vccd1 vccd1
+ _14376_/D sky130_fd_sc_hd__o221a_1
XFILLER_182_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _13547_/Q _09048_/X _08970_/X _09049_/X _09045_/X vssd1 vssd1 vccd1 vccd1
+ _13547_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08001_ _14066_/Q _07999_/X _07771_/X _08000_/X _07995_/X vssd1 vssd1 vccd1 vccd1
+ _14066_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09952_ _09952_/A vssd1 vssd1 vccd1 vccd1 _09952_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08903_ _13612_/Q _08894_/X _08829_/X _08897_/X _08900_/X vssd1 vssd1 vccd1 vccd1
+ _13612_/D sky130_fd_sc_hd__o221a_1
XFILLER_48_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09883_ _09883_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__or2_2
XFILLER_44_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08834_ _08877_/A vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _13686_/Q _08758_/X _08508_/X _08760_/X _08761_/X vssd1 vssd1 vccd1 vccd1
+ _13686_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07716_ _14204_/Q _07704_/X _07714_/X _07706_/X _07715_/X vssd1 vssd1 vccd1 vccd1
+ _14204_/D sky130_fd_sc_hd__o221a_1
XPHY_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _08728_/A vssd1 vssd1 vccd1 vccd1 _08696_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07647_ _14242_/Q _07644_/X _07323_/X _07646_/X _07640_/X vssd1 vssd1 vccd1 vccd1
+ _14242_/D sky130_fd_sc_hd__o221a_1
XPHY_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ _14278_/Q _07571_/X _07330_/X _07573_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _14278_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _13397_/Q _09310_/X _08158_/A _09311_/X _09314_/X vssd1 vssd1 vccd1 vccd1
+ _13397_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06529_ _06823_/A vssd1 vssd1 vccd1 vccd1 _06530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _13436_/Q _09241_/X _08954_/X _09242_/X _09244_/X vssd1 vssd1 vccd1 vccd1
+ _13436_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09179_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11210_ _13598_/Q vssd1 vssd1 vccd1 vccd1 _11210_/Y sky130_fd_sc_hd__inv_2
X_12190_ vssd1 vssd1 vccd1 vccd1 _12190_/HI _12190_/LO sky130_fd_sc_hd__conb_1
XFILLER_159_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _14345_/Q vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11072_ _13478_/Q vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput100 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _07086_/B sky130_fd_sc_hd__buf_4
XPHY_7121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput111 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__buf_4
XFILLER_27_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _13380_/Q _10023_/B vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__nand2_1
Xinput122 la_data_in[5] vssd1 vssd1 vccd1 vccd1 _07803_/A sky130_fd_sc_hd__buf_6
XFILLER_46_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 la_data_in[6] vssd1 vssd1 vccd1 vccd1 _08989_/D sky130_fd_sc_hd__buf_6
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput144 la_data_in[7] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__buf_1
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 la_data_in[8] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__buf_1
XPHY_7176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 la_data_in[9] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_1
XPHY_7187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 la_oenb[109] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__buf_1
XFILLER_40_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 la_oenb[119] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__buf_1
XPHY_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 la_oenb[13] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__buf_1
XFILLER_40_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11974_ _11972_/Y _10220_/A _11973_/Y _10223_/A vssd1 vssd1 vccd1 vccd1 _11974_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _14146_/CLK _13713_/D vssd1 vssd1 vccd1 vccd1 _13713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10925_ _11399_/A vssd1 vssd1 vccd1 vccd1 _10925_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13644_ _14143_/CLK _13644_/D vssd1 vssd1 vccd1 vccd1 _13644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10856_ _13513_/Q vssd1 vssd1 vccd1 vccd1 _10856_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13575_ _14130_/CLK _13575_/D vssd1 vssd1 vccd1 vccd1 _13575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ _14259_/Q vssd1 vssd1 vccd1 vccd1 _10787_/Y sky130_fd_sc_hd__inv_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12526_ _13374_/Q _10037_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12457_ _12456_/X _06927_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12457_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ _11408_/A vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__clkbuf_2
Xoutput607 _13264_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_2
X_12388_ _12387_/X _13209_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14127_ _14130_/CLK _14127_/D vssd1 vssd1 vccd1 vccd1 _14127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11339_ _11337_/Y _11203_/X _11338_/Y _11205_/X vssd1 vssd1 vccd1 vccd1 _11339_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ _14139_/CLK _14058_/D vssd1 vssd1 vccd1 vccd1 _14058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13009_ _12584_/X _13008_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06880_ _06956_/A vssd1 vssd1 vccd1 vccd1 _06880_/X sky130_fd_sc_hd__buf_1
XFILLER_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08550_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07501_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08481_ _13819_/Q _08415_/A _08268_/X _08417_/A _08480_/X vssd1 vssd1 vccd1 vccd1
+ _13819_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07432_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07363_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07363_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _13519_/Q _09095_/X _08942_/X _09096_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _13519_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07294_ _14410_/Q _07290_/X _06831_/X _07291_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _14410_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09033_ _13556_/Q _09030_/X _08948_/X _09031_/X _09027_/X vssd1 vssd1 vccd1 vccd1
+ _13556_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09935_ _09899_/A _09899_/B _09934_/Y vssd1 vssd1 vccd1 vccd1 _09935_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09866_ _13302_/Q vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__inv_2
XFILLER_63_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08817_ _08876_/A vssd1 vssd1 vccd1 vccd1 _08818_/A sky130_fd_sc_hd__clkbuf_2
XPHY_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09797_ _13344_/Q vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__inv_2
XPHY_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08748_/A vssd1 vssd1 vccd1 vccd1 _08748_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _13273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08679_ _08679_/A vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _14102_/Q vssd1 vssd1 vccd1 vccd1 _10710_/Y sky130_fd_sc_hd__inv_2
XPHY_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11690_ _14161_/Q vssd1 vssd1 vccd1 vccd1 _11690_/Y sky130_fd_sc_hd__inv_2
XPHY_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _10639_/Y _10512_/X _10640_/Y _10515_/X vssd1 vssd1 vccd1 vccd1 _10641_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13360_ _14639_/CLK _13360_/D vssd1 vssd1 vccd1 vccd1 _13360_/Q sky130_fd_sc_hd__dfxtp_1
X_10572_ _13748_/Q vssd1 vssd1 vccd1 vccd1 _10572_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _10797_/Y _14532_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__mux2_2
XFILLER_52_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _13877_/CLK _13291_/D vssd1 vssd1 vccd1 vccd1 _13291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12242_ _12242_/A vssd1 vssd1 vccd1 vccd1 _12242_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12173_ vssd1 vssd1 vccd1 vccd1 _12173_/HI _12173_/LO sky130_fd_sc_hd__conb_1
XFILLER_155_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _11119_/Y _10923_/X _11120_/Y _10925_/X _11123_/X vssd1 vssd1 vccd1 vccd1
+ _11159_/A sky130_fd_sc_hd__o221a_1
XFILLER_155_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11055_ _11045_/Y _10940_/X _11048_/X _11051_/X _11054_/X vssd1 vssd1 vccd1 vccd1
+ _11077_/C sky130_fd_sc_hd__o2111a_4
XFILLER_190_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10006_ _13374_/Q _10006_/B vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _13973_/Q vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__inv_2
XPHY_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _14301_/Q vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__inv_2
XPHY_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11888_ _14517_/Q vssd1 vssd1 vccd1 vccd1 _11888_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13627_ _14119_/CLK _13627_/D vssd1 vssd1 vccd1 vccd1 _13627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10839_ _10839_/A _10839_/B _10839_/C _10839_/D vssd1 vssd1 vccd1 vccd1 _10839_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_109_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ _14114_/CLK _13558_/D vssd1 vssd1 vccd1 vccd1 _13558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12509_ _12508_/X _10058_/Y _12509_/S vssd1 vssd1 vccd1 vccd1 _12509_/X sky130_fd_sc_hd__mux2_8
XFILLER_172_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13489_ _14470_/CLK _13489_/D vssd1 vssd1 vccd1 vccd1 _13489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput404 _12204_/X vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__clkbuf_2
Xoutput415 _12094_/LO vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput426 _12242_/A vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput437 _12079_/LO vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput448 _12235_/X vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput459 _12245_/X vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07981_ _14077_/Q _07974_/X _07742_/X _07975_/X _07978_/X vssd1 vssd1 vccd1 vccd1
+ _14077_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09720_ _09718_/X _09719_/X _09718_/X _09719_/X vssd1 vssd1 vccd1 vccd1 _09720_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06932_ _06935_/A _06932_/B vssd1 vssd1 vccd1 vccd1 _14580_/D sky130_fd_sc_hd__nor2_1
XFILLER_60_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09651_ _06875_/Y _14562_/Q _14594_/Q _06996_/Y vssd1 vssd1 vccd1 vccd1 _09651_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06863_ _06877_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _14598_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08602_ _08645_/A vssd1 vssd1 vccd1 vccd1 _08637_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _09586_/A _12328_/X vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__and2_1
XFILLER_97_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06794_ _14616_/Q _06787_/X _06793_/X _06790_/X _06785_/X vssd1 vssd1 vccd1 vccd1
+ _14616_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ _13801_/Q _08526_/X _08532_/X _08528_/X _08524_/X vssd1 vssd1 vccd1 vccd1
+ _13801_/D sky130_fd_sc_hd__o221a_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08464_ _13830_/Q _08460_/X _08167_/X _08461_/X _08457_/X vssd1 vssd1 vccd1 vccd1
+ _13830_/D sky130_fd_sc_hd__o221a_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07415_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07415_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ _13867_/Q _08388_/X _08171_/X _08389_/X _08392_/X vssd1 vssd1 vccd1 vccd1
+ _13867_/D sky130_fd_sc_hd__o221a_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07346_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07346_/X sky130_fd_sc_hd__buf_2
XFILLER_71_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07277_ _14421_/Q _07274_/X _06793_/X _07275_/X _07271_/X vssd1 vssd1 vccd1 vccd1
+ _14421_/D sky130_fd_sc_hd__o221a_1
XFILLER_203_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09016_ _13567_/Q _09014_/X _08917_/X _09015_/X _09011_/X vssd1 vssd1 vccd1 vccd1
+ _13567_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09918_ _13315_/Q vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__inv_2
XFILLER_82_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _09771_/A _09771_/B _09772_/B vssd1 vssd1 vccd1 vccd1 _09849_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_41_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12860_ _12526_/X input345/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11811_ _13611_/Q vssd1 vssd1 vccd1 vccd1 _11811_/Y sky130_fd_sc_hd__inv_2
XPHY_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _09533_/X _12790_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13216_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14611_/CLK _14530_/D vssd1 vssd1 vccd1 vccd1 _14530_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _13454_/Q vssd1 vssd1 vccd1 vccd1 _11742_/Y sky130_fd_sc_hd__inv_2
XPHY_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14595_/CLK _14461_/D vssd1 vssd1 vccd1 vccd1 _14461_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11673_ _11673_/A vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13412_ _14178_/CLK _13412_/D vssd1 vssd1 vccd1 vccd1 _13412_/Q sky130_fd_sc_hd__dfxtp_1
X_10624_ _13199_/Q _10539_/X _14022_/Q _10469_/X _10623_/X vssd1 vssd1 vccd1 vccd1
+ _10624_/X sky130_fd_sc_hd__a221o_4
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14392_ _14629_/CLK _14392_/D vssd1 vssd1 vccd1 vccd1 _14392_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343_ _14538_/CLK _13343_/D vssd1 vssd1 vccd1 vccd1 _13343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ _14137_/Q vssd1 vssd1 vccd1 vccd1 _10555_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13274_ _13371_/CLK _13274_/D vssd1 vssd1 vccd1 vccd1 _13274_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10486_ _11675_/A vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__buf_2
XFILLER_182_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12225_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12156_ vssd1 vssd1 vccd1 vccd1 _12156_/HI _12156_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11107_ _14188_/Q vssd1 vssd1 vccd1 vccd1 _11107_/Y sky130_fd_sc_hd__inv_2
X_12087_ vssd1 vssd1 vccd1 vccd1 _12087_/HI _12087_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11038_ _13673_/Q vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989_ _12574_/X _12988_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__mux2_1
XPHY_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07200_ _14462_/Q _07193_/X _06784_/X _07194_/X _07197_/X vssd1 vssd1 vccd1 vccd1
+ _14462_/D sky130_fd_sc_hd__o221a_1
X_08180_ _13981_/Q _08174_/X _08179_/X _08176_/X _08172_/X vssd1 vssd1 vccd1 vccd1
+ _13981_/D sky130_fd_sc_hd__o221a_1
XFILLER_158_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07131_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07131_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07062_ _07062_/A vssd1 vssd1 vccd1 vccd1 _07062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07964_ _08007_/A vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__buf_6
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09701_/Y _09702_/X _09701_/Y _09702_/X vssd1 vssd1 vccd1 vccd1 _09703_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06915_ _14584_/Q vssd1 vssd1 vccd1 vccd1 _06915_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07895_ _14125_/Q _07892_/X _07719_/X _07894_/X _07886_/X vssd1 vssd1 vccd1 vccd1
+ _14125_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09634_ _09632_/X _09633_/X _09632_/X _09633_/X vssd1 vssd1 vccd1 vccd1 _09634_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06846_ _14601_/Q _06530_/A _06845_/X _06532_/A _06838_/X vssd1 vssd1 vccd1 vccd1
+ _14601_/D sky130_fd_sc_hd__o221a_1
XFILLER_186_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09565_ _09573_/A _12355_/X vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__and2_1
X_06777_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08142_/A sky130_fd_sc_hd__buf_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _13808_/Q _08513_/X _08514_/X _08515_/X _08511_/X vssd1 vssd1 vccd1 vccd1
+ _13808_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _13265_/Q _09493_/X _12260_/X _09494_/X vssd1 vssd1 vccd1 vccd1 _13265_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _13841_/Q _08444_/X _08140_/X _08445_/X _08441_/X vssd1 vssd1 vccd1 vccd1
+ _13841_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _13877_/Q _08371_/X _08146_/X _08372_/X _08375_/X vssd1 vssd1 vccd1 vccd1
+ _13877_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07329_ _14396_/Q _07322_/X _07031_/X _07325_/X _07319_/X vssd1 vssd1 vccd1 vccd1
+ _14396_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10340_ _10340_/A _10340_/B _10340_/C _10340_/D vssd1 vssd1 vccd1 vccd1 _10340_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_137_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10271_ _13976_/Q vssd1 vssd1 vccd1 vccd1 _10271_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12010_ _13733_/Q _10173_/A _14052_/Q _10203_/A _12009_/X vssd1 vssd1 vccd1 vccd1
+ _12010_/X sky130_fd_sc_hd__a221o_2
XFILLER_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13961_ _14110_/CLK _13961_/D vssd1 vssd1 vccd1 vccd1 _13961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12912_ _12539_/X input348/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13892_ _14130_/CLK _13892_/D vssd1 vssd1 vccd1 vccd1 _13892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12843_ _12521_/X _12842_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12774_ _09522_/X _12773_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12774_/X sky130_fd_sc_hd__mux2_1
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14513_ _14629_/CLK _14513_/D vssd1 vssd1 vccd1 vccd1 _14513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11725_ _11723_/Y _11673_/X _11724_/Y _11675_/X vssd1 vssd1 vccd1 vccd1 _11725_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _14481_/CLK _14444_/D vssd1 vssd1 vccd1 vccd1 _14444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11652_/Y _11653_/X _11654_/Y _11655_/X vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _13625_/Q vssd1 vssd1 vccd1 vccd1 _10607_/Y sky130_fd_sc_hd__inv_2
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14375_ _14627_/CLK _14375_/D vssd1 vssd1 vccd1 vccd1 _14375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11587_ _11585_/Y _11459_/X _11586_/Y _11461_/X vssd1 vssd1 vccd1 vccd1 _11587_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _13877_/CLK _13326_/D vssd1 vssd1 vccd1 vccd1 _13326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10538_ _10528_/Y _10445_/X _10531_/X _10534_/X _10537_/X vssd1 vssd1 vccd1 vccd1
+ _10561_/C sky130_fd_sc_hd__o2111a_4
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13257_ _14639_/CLK _13257_/D vssd1 vssd1 vccd1 vccd1 _13257_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_48_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10469_ _11429_/A vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12208_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13188_ _13185_/X _12507_/X _13186_/X _13187_/X _12510_/S _10058_/B vssd1 vssd1 vccd1
+ vccd1 _13188_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12139_ vssd1 vssd1 vccd1 vccd1 _12139_/HI _12139_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater704 _12853_/S vssd1 vssd1 vccd1 vccd1 _13113_/S sky130_fd_sc_hd__buf_8
XFILLER_26_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06700_ _06699_/Y _06646_/X _06699_/Y _06646_/X vssd1 vssd1 vccd1 vccd1 _06700_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07680_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07680_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06631_ _06624_/X _06630_/X _06624_/X _06630_/X vssd1 vssd1 vccd1 vccd1 _06632_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _09351_/A _12863_/X vssd1 vssd1 vccd1 vccd1 _13374_/D sky130_fd_sc_hd__and2_1
X_06562_ _06562_/A vssd1 vssd1 vccd1 vccd1 _06562_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08301_ _13921_/Q _08293_/X _08132_/X _08294_/X _08297_/X vssd1 vssd1 vccd1 vccd1
+ _13921_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _13419_/Q _09275_/X _07710_/A _09277_/X _09280_/X vssd1 vssd1 vccd1 vccd1
+ _13419_/D sky130_fd_sc_hd__o221a_1
X_06493_ _06493_/A _06493_/B _06493_/C _06493_/D vssd1 vssd1 vccd1 vccd1 _06499_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08232_ _13959_/Q _08229_/X _08137_/X _08230_/X _08231_/X vssd1 vssd1 vccd1 vccd1
+ _13959_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08163_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07114_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07114_/X sky130_fd_sc_hd__buf_2
X_08094_ _08174_/A vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ _07062_/A vssd1 vssd1 vccd1 vccd1 _07045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _13577_/Q _08993_/X _08895_/X _08995_/X _08986_/X vssd1 vssd1 vccd1 vccd1
+ _13577_/D sky130_fd_sc_hd__o221a_1
XFILLER_125_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _14094_/Q _07882_/A _07798_/X _07884_/A _07946_/X vssd1 vssd1 vccd1 vccd1
+ _14094_/D sky130_fd_sc_hd__o221a_1
XPHY_6838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07878_ _08814_/A _07878_/B _09271_/C _08091_/D vssd1 vssd1 vccd1 vccd1 _11655_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_95_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09617_ _06924_/Y _06989_/X _14582_/Q _14564_/Q vssd1 vssd1 vccd1 vccd1 _09617_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06829_ _06853_/A _06829_/B vssd1 vssd1 vccd1 vccd1 _06829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09548_ _09544_/X _09547_/X _13275_/Q _09545_/X vssd1 vssd1 vccd1 vccd1 _13243_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09479_ _09479_/A vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__clkbuf_2
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _13683_/Q vssd1 vssd1 vccd1 vccd1 _11510_/Y sky130_fd_sc_hd__inv_2
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12490_ _12489_/X _06970_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12490_/X sky130_fd_sc_hd__mux2_2
XFILLER_12_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _11441_/A vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14160_ _14291_/CLK _14160_/D vssd1 vssd1 vccd1 vccd1 _14160_/Q sky130_fd_sc_hd__dfxtp_1
X_11372_ _11370_/Y _11188_/X _11371_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11372_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _12633_/X _13110_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13111_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10323_ _14601_/Q vssd1 vssd1 vccd1 vccd1 _10323_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14091_ _14169_/CLK _14091_/D vssd1 vssd1 vccd1 vccd1 _14091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _13041_/X _12600_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10254_ _10211_/X _10254_/B _10254_/C _10254_/D vssd1 vssd1 vccd1 vccd1 _10255_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10185_ _10179_/Y _10181_/X _10182_/Y _10184_/X vssd1 vssd1 vccd1 vccd1 _10185_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13944_ _14100_/CLK _13944_/D vssd1 vssd1 vccd1 vccd1 _13944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13875_ _13877_/CLK _13875_/D vssd1 vssd1 vccd1 vccd1 _13875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12826_ _10048_/X _12825_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12826_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12757_ _09554_/X _12756_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11708_ _13967_/Q vssd1 vssd1 vccd1 vccd1 _11708_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ _09593_/X input352/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14427_ _14595_/CLK _14427_/D vssd1 vssd1 vccd1 vccd1 _14427_/Q sky130_fd_sc_hd__dfxtp_1
X_11639_ _11639_/A vssd1 vssd1 vccd1 vccd1 _11639_/X sky130_fd_sc_hd__buf_2
XFILLER_200_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14358_ _14629_/CLK _14358_/D vssd1 vssd1 vccd1 vccd1 _14358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13309_ _14538_/CLK _13309_/D vssd1 vssd1 vccd1 vccd1 _13309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14289_ _14325_/CLK _14289_/D vssd1 vssd1 vccd1 vccd1 _14289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ _13642_/Q _08844_/X _08521_/X _08845_/X _08847_/X vssd1 vssd1 vccd1 vccd1
+ _13642_/D sky130_fd_sc_hd__o221a_1
XFILLER_170_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07801_ _14171_/Q _07704_/A _07800_/X _07706_/A _07794_/X vssd1 vssd1 vccd1 vccd1
+ _14171_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08781_ _13676_/Q _08775_/X _08534_/X _08776_/X _08777_/X vssd1 vssd1 vccd1 vccd1
+ _13676_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07732_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07732_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07663_ _14232_/Q _07661_/X _07349_/X _07662_/X _07658_/X vssd1 vssd1 vccd1 vccd1
+ _14232_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06614_ _06614_/A vssd1 vssd1 vccd1 vccd1 _06614_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07594_ _14269_/Q _07589_/X _07354_/X _07590_/X _07593_/X vssd1 vssd1 vccd1 vccd1
+ _14269_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09333_ _13387_/Q _09326_/X _08183_/A _09327_/X _09330_/X vssd1 vssd1 vccd1 vccd1
+ _13387_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06545_ _06545_/A vssd1 vssd1 vccd1 vccd1 _06545_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09264_ _13426_/Q _09257_/X _08979_/X _09258_/X _09260_/X vssd1 vssd1 vccd1 vccd1
+ _13426_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08215_ _13969_/Q _08211_/X _08110_/X _08213_/X _08214_/X vssd1 vssd1 vccd1 vccd1
+ _13969_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09195_ _13465_/Q _09188_/X _08979_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1
+ _13465_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ _08146_/A vssd1 vssd1 vccd1 vccd1 _08146_/X sky130_fd_sc_hd__buf_4
XFILLER_147_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08077_ _14023_/Q _08069_/X _07780_/X _08070_/X _08075_/X vssd1 vssd1 vccd1 vccd1
+ _14023_/D sky130_fd_sc_hd__o221a_1
XFILLER_49_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07028_ _07028_/A vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput304 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _06493_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput315 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _06494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput326 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _06507_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput337 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input337/X sky130_fd_sc_hd__clkbuf_4
XPHY_7358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__buf_4
Xinput348 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 input348/X sky130_fd_sc_hd__buf_6
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput359 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input359/X sky130_fd_sc_hd__clkbuf_4
XPHY_6635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _14091_/Q vssd1 vssd1 vccd1 vccd1 _11990_/Y sky130_fd_sc_hd__inv_2
XPHY_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10941_ _13756_/Q vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__inv_2
XPHY_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13660_ _14047_/CLK _13660_/D vssd1 vssd1 vccd1 vccd1 _13660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10872_ _10867_/Y _10735_/X _10868_/Y _10737_/X _10871_/X vssd1 vssd1 vccd1 vccd1
+ _10879_/C sky130_fd_sc_hd__o221a_1
XFILLER_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _09852_/X _13323_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _14188_/CLK _13591_/D vssd1 vssd1 vccd1 vccd1 _13591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12542_ _09964_/Y _13294_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12473_ _12509_/X _06952_/Y _12473_/S vssd1 vssd1 vccd1 vccd1 _12473_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14212_ _14325_/CLK _14212_/D vssd1 vssd1 vccd1 vccd1 _14212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11424_ _11424_/A vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 _12304_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14143_/CLK _14143_/D vssd1 vssd1 vccd1 vccd1 _14143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11355_ _14077_/Q vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10306_ _13385_/Q _10305_/X _13697_/Q _10173_/X vssd1 vssd1 vccd1 vccd1 _10306_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14074_ _14459_/CLK _14074_/D vssd1 vssd1 vccd1 vccd1 _14074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11286_ _14114_/Q vssd1 vssd1 vccd1 vccd1 _11286_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13025_ _12592_/X _13024_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _13025_/X sky130_fd_sc_hd__mux2_1
X_10237_ _10237_/A vssd1 vssd1 vccd1 vccd1 _10237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _10168_/A vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__inv_2
XFILLER_187_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10099_ _10099_/A _10138_/A vssd1 vssd1 vccd1 vccd1 _12473_/S sky130_fd_sc_hd__or2_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13927_ _14139_/CLK _13927_/D vssd1 vssd1 vccd1 vccd1 _13927_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13858_ _14095_/CLK _13858_/D vssd1 vssd1 vccd1 vccd1 _13858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _12514_/X _12808_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13789_ _14120_/CLK _13789_/D vssd1 vssd1 vccd1 vccd1 _13789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _08000_/A vssd1 vssd1 vccd1 vccd1 _08000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09951_ _13300_/Q _09949_/Y _09895_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ _13613_/Q _08894_/X _08827_/X _08897_/X _08900_/X vssd1 vssd1 vccd1 vccd1
+ _13613_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09882_ _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__or2_2
XFILLER_48_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ _08833_/A vssd1 vssd1 vccd1 vccd1 _08833_/X sky130_fd_sc_hd__buf_4
XFILLER_83_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08764_ _13687_/Q _08758_/X _08606_/X _08760_/X _08761_/X vssd1 vssd1 vccd1 vccd1
+ _13687_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07715_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07715_/X sky130_fd_sc_hd__buf_2
XPHY_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08695_ _08879_/A vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07646_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07646_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07577_ _14279_/Q _07571_/X _07428_/X _07573_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _14279_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09316_ _13398_/Q _09310_/X _09035_/X _09311_/X _09314_/X vssd1 vssd1 vccd1 vccd1
+ _13398_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06528_ _06811_/A vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__inv_2
XFILLER_146_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09247_ _13437_/Q _09241_/X _09035_/X _09242_/X _09244_/X vssd1 vssd1 vccd1 vccd1
+ _13437_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _13475_/Q _09171_/X _08954_/X _09172_/X _09173_/X vssd1 vssd1 vccd1 vccd1
+ _13475_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ _14001_/Q _08122_/X _08128_/X _08124_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _14001_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11140_ _14501_/Q vssd1 vssd1 vccd1 vccd1 _11140_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11071_ _14148_/Q vssd1 vssd1 vccd1 vccd1 _11071_/Y sky130_fd_sc_hd__inv_2
XPHY_7100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput101 la_data_in[40] vssd1 vssd1 vccd1 vccd1 _06559_/A sky130_fd_sc_hd__buf_2
XFILLER_81_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10022_ _10022_/A vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__inv_2
Xinput112 la_data_in[50] vssd1 vssd1 vccd1 vccd1 _06639_/A sky130_fd_sc_hd__buf_2
XPHY_7133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput123 la_data_in[60] vssd1 vssd1 vccd1 vccd1 _06546_/A sky130_fd_sc_hd__buf_2
XFILLER_27_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput134 la_data_in[70] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__buf_1
XFILLER_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 la_data_in[80] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__buf_1
XPHY_7166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 la_data_in[90] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__buf_1
XFILLER_44_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput167 la_oenb[0] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__buf_1
XPHY_7188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput178 la_oenb[10] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__buf_1
XPHY_7199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 la_oenb[11] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_hd__buf_1
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ _14402_/Q vssd1 vssd1 vccd1 vccd1 _11973_/Y sky130_fd_sc_hd__inv_2
XPHY_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _14146_/CLK _13712_/D vssd1 vssd1 vccd1 vccd1 _13712_/Q sky130_fd_sc_hd__dfxtp_1
X_10924_ _13437_/Q vssd1 vssd1 vccd1 vccd1 _10924_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13643_ _14143_/CLK _13643_/D vssd1 vssd1 vccd1 vccd1 _13643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10855_ _13988_/Q vssd1 vssd1 vccd1 vccd1 _10855_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13574_ _14130_/CLK _13574_/D vssd1 vssd1 vccd1 vccd1 _13574_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _14181_/Q vssd1 vssd1 vccd1 vccd1 _10786_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12525_ _13359_/Q _10038_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ _12455_/X _06927_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__mux2_1
X_11407_ _11407_/A vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12387_ _13209_/Q _12386_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14126_ _14130_/CLK _14126_/D vssd1 vssd1 vccd1 vccd1 _14126_/Q sky130_fd_sc_hd__dfxtp_1
X_11338_ _14388_/Q vssd1 vssd1 vccd1 vccd1 _11338_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ _14139_/CLK _14057_/D vssd1 vssd1 vccd1 vccd1 _14057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11269_ _11264_/Y _11219_/X _11265_/Y _11221_/X _11268_/X vssd1 vssd1 vccd1 vccd1
+ _11270_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13008_ _12584_/X input339/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07500_ _07542_/A vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__buf_4
XFILLER_110_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08480_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08480_/X sky130_fd_sc_hd__buf_2
XFILLER_36_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07431_ _14355_/Q _07422_/X _07332_/X _07424_/X _07425_/X vssd1 vssd1 vccd1 vccd1
+ _14355_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07362_ _08150_/A vssd1 vssd1 vccd1 vccd1 _07362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09101_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07293_ _14411_/Q _07290_/X _07073_/X _07291_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _14411_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09032_ _13557_/Q _09030_/X _08945_/X _09031_/X _09027_/X vssd1 vssd1 vccd1 vccd1
+ _13557_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _09934_/A vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09865_ _13303_/Q vssd1 vssd1 vccd1 vccd1 _09897_/A sky130_fd_sc_hd__inv_2
XFILLER_24_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08816_ _08877_/A vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__inv_2
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09796_ _09847_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09796_/X sky130_fd_sc_hd__and2_4
XPHY_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08747_ _08800_/A vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__clkbuf_2
XPHY_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _13256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08678_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08679_/A sky130_fd_sc_hd__buf_2
XPHY_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07629_ _09131_/A vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _14451_/Q vssd1 vssd1 vccd1 vccd1 _10640_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10571_ _13943_/Q vssd1 vssd1 vccd1 vccd1 _10571_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12310_ _10839_/Y _14533_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12310_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13290_ _13877_/CLK _13290_/D vssd1 vssd1 vccd1 vccd1 _13290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12241_ _12241_/A vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12172_ vssd1 vssd1 vccd1 vccd1 _12172_/HI _12172_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11123_ _11121_/Y _10927_/X _11122_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _11123_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_190_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11054_ _11052_/Y _10952_/X _11053_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _11054_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10005_ _10005_/A vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__inv_2
XFILLER_209_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11956_ _13420_/Q _11747_/A _13739_/Q _09601_/A _11955_/X vssd1 vssd1 vccd1 vccd1
+ _11989_/B sky130_fd_sc_hd__a221oi_2
XPHY_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ _10902_/Y _10725_/X _10903_/Y _10727_/X _10906_/X vssd1 vssd1 vccd1 vccd1
+ _10920_/B sky130_fd_sc_hd__o221a_4
X_11887_ _13730_/Q _10173_/A _14049_/Q _10203_/A _11886_/X vssd1 vssd1 vccd1 vccd1
+ _11887_/X sky130_fd_sc_hd__a221o_4
XFILLER_33_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13626_ _14119_/CLK _13626_/D vssd1 vssd1 vccd1 vccd1 _13626_/Q sky130_fd_sc_hd__dfxtp_1
X_10838_ _10819_/X _10838_/B _10838_/C _10838_/D vssd1 vssd1 vccd1 vccd1 _10839_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_92_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10769_ _14103_/Q vssd1 vssd1 vccd1 vccd1 _10769_/Y sky130_fd_sc_hd__inv_2
X_13557_ _14114_/CLK _13557_/D vssd1 vssd1 vccd1 vccd1 _13557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12508_ _13184_/X _13188_/X _12508_/S vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__mux2_1
X_13488_ _14470_/CLK _13488_/D vssd1 vssd1 vccd1 vccd1 _13488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12439_ _12438_/X _06906_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12439_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput405 _12205_/X vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput416 _12095_/LO vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput427 _12243_/A vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput438 _12080_/LO vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput449 _12236_/X vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14109_ _14110_/CLK _14109_/D vssd1 vssd1 vccd1 vccd1 _14109_/Q sky130_fd_sc_hd__dfxtp_1
X_07980_ _14078_/Q _07974_/X _07740_/X _07975_/X _07978_/X vssd1 vssd1 vccd1 vccd1
+ _14078_/D sky130_fd_sc_hd__o221a_1
XFILLER_64_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06931_ _06919_/X _12302_/X _06930_/Y _06921_/X vssd1 vssd1 vccd1 vccd1 _06932_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09650_ _09650_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _12486_/S sky130_fd_sc_hd__nand2_4
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06862_ _06857_/X _12284_/X _06858_/Y _06861_/X vssd1 vssd1 vccd1 vccd1 _06863_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08601_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08601_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09581_ _09570_/X _09580_/X _13262_/Q _09571_/X vssd1 vssd1 vccd1 vccd1 _13230_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06793_ _08153_/A vssd1 vssd1 vccd1 vccd1 _06793_/X sky130_fd_sc_hd__buf_4
XFILLER_209_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08532_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08532_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08463_ _13831_/Q _08460_/X _08165_/X _08461_/X _08457_/X vssd1 vssd1 vccd1 vccd1
+ _13831_/D sky130_fd_sc_hd__o221a_1
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07414_ _07414_/A vssd1 vssd1 vccd1 vccd1 _07414_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08394_ _13868_/Q _08388_/X _08169_/X _08389_/X _08392_/X vssd1 vssd1 vccd1 vccd1
+ _13868_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07345_ _08132_/A vssd1 vssd1 vccd1 vccd1 _07345_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07276_ _14422_/Q _07274_/X _06789_/X _07275_/X _07271_/X vssd1 vssd1 vccd1 vccd1
+ _14422_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09015_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ _13314_/Q _09913_/Y _09919_/B vssd1 vssd1 vccd1 vccd1 _09917_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09848_ _13320_/Q _13319_/Q _09771_/B vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__or2_1
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11810_ _14320_/Q vssd1 vssd1 vccd1 vccd1 _11810_/Y sky130_fd_sc_hd__inv_2
XPHY_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12790_ _09533_/X _12789_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _14085_/Q vssd1 vssd1 vccd1 vccd1 _11741_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _14629_/Q vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14460_ _14595_/CLK _14460_/D vssd1 vssd1 vccd1 vccd1 _14460_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _13547_/Q _10471_/X _13788_/Q _10473_/X vssd1 vssd1 vccd1 vccd1 _10623_/X
+ sky130_fd_sc_hd__a22o_1
X_13411_ _14183_/CLK _13411_/D vssd1 vssd1 vccd1 vccd1 _13411_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _14629_/CLK _14391_/D vssd1 vssd1 vccd1 vccd1 _14391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _14538_/CLK _13342_/D vssd1 vssd1 vccd1 vccd1 _13342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10554_ _13903_/Q vssd1 vssd1 vccd1 vccd1 _10554_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13273_ _13368_/CLK _13273_/D vssd1 vssd1 vccd1 vccd1 _13273_/Q sky130_fd_sc_hd__dfxtp_4
X_10485_ _14370_/Q vssd1 vssd1 vccd1 vccd1 _10485_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12224_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ vssd1 vssd1 vccd1 vccd1 _12155_/HI _12155_/LO sky130_fd_sc_hd__conb_1
XFILLER_194_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11106_ _13596_/Q vssd1 vssd1 vccd1 vccd1 _11106_/Y sky130_fd_sc_hd__inv_2
X_12086_ vssd1 vssd1 vccd1 vccd1 _12086_/HI _12086_/LO sky130_fd_sc_hd__conb_1
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11037_ _13439_/Q vssd1 vssd1 vccd1 vccd1 _11037_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12988_ _12574_/X input345/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11939_ _11937_/Y _10234_/A _11938_/Y _10237_/A vssd1 vssd1 vccd1 vccd1 _11939_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_206_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13609_ _14481_/CLK _13609_/D vssd1 vssd1 vccd1 vccd1 _13609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14589_ _14621_/CLK _14589_/D vssd1 vssd1 vccd1 vccd1 _14589_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _07130_/A vssd1 vssd1 vccd1 vccd1 _07169_/A sky130_fd_sc_hd__buf_2
XFILLER_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07061_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _14087_/Q _07955_/X _07714_/X _07957_/X _07960_/X vssd1 vssd1 vccd1 vccd1
+ _14087_/D sky130_fd_sc_hd__o221a_1
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ _06906_/Y _14583_/Q _14587_/Q _06920_/Y vssd1 vssd1 vccd1 vccd1 _09702_/X
+ sky130_fd_sc_hd__o22a_1
X_06914_ _06917_/A _06914_/B vssd1 vssd1 vccd1 vccd1 _14585_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07894_ _07927_/A vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06845_ _08188_/A vssd1 vssd1 vccd1 vccd1 _06845_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _06999_/Y _10057_/A _14561_/Q _14560_/Q vssd1 vssd1 vccd1 vccd1 _09633_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09564_ _09557_/X _09563_/X _13269_/Q _09558_/X vssd1 vssd1 vccd1 vccd1 _13237_/D
+ sky130_fd_sc_hd__o22a_1
X_06776_ _14621_/Q _06769_/X _06775_/X _06772_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _14621_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08515_ _08554_/A vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09495_ _13266_/Q _09493_/X _12261_/X _09494_/X vssd1 vssd1 vccd1 vccd1 _13266_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08446_ _13842_/Q _08444_/X _08137_/X _08445_/X _08441_/X vssd1 vssd1 vccd1 vccd1
+ _13842_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ _13878_/Q _08371_/X _08144_/X _08372_/X _08375_/X vssd1 vssd1 vccd1 vccd1
+ _13878_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07328_ _14397_/Q _07322_/X _07327_/X _07325_/X _07319_/X vssd1 vssd1 vccd1 vccd1
+ _14397_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07259_ _14432_/Q _07257_/X _06753_/X _07258_/X _07254_/X vssd1 vssd1 vccd1 vccd1
+ _14432_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ _10268_/Y _10188_/X _10269_/Y _10191_/X vssd1 vssd1 vccd1 vccd1 _10270_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13960_ _14110_/CLK _13960_/D vssd1 vssd1 vccd1 vccd1 _13960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12911_ _12538_/X _12910_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13891_ _14100_/CLK _13891_/D vssd1 vssd1 vccd1 vccd1 _13891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12842_ _12521_/X _12841_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12773_ _09522_/X _12772_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14629_/CLK _14512_/D vssd1 vssd1 vccd1 vccd1 _14512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11724_ _14396_/Q vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14443_ _14481_/CLK _14443_/D vssd1 vssd1 vccd1 vccd1 _14443_/Q sky130_fd_sc_hd__dfxtp_1
X_11655_ _11655_/A vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10606_ _13664_/Q vssd1 vssd1 vccd1 vccd1 _10606_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11586_ _14471_/Q vssd1 vssd1 vccd1 vccd1 _11586_/Y sky130_fd_sc_hd__inv_2
X_14374_ _14627_/CLK _14374_/D vssd1 vssd1 vccd1 vccd1 _14374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10537_ _10535_/Y _10462_/X _10536_/Y _10465_/X vssd1 vssd1 vccd1 vccd1 _10537_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13325_ _13877_/CLK _13325_/D vssd1 vssd1 vccd1 vccd1 _13325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10468_ _11663_/A vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__clkbuf_2
X_13256_ _13352_/CLK _13256_/D vssd1 vssd1 vccd1 vccd1 _13256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_48_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13187_ _14569_/Q _14570_/Q _14567_/Q _14568_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13187_/X sky130_fd_sc_hd__mux4_2
XFILLER_151_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10399_ _10397_/Y _10195_/X _10398_/Y _10198_/X vssd1 vssd1 vccd1 vccd1 _10399_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12138_ vssd1 vssd1 vccd1 vccd1 _12138_/HI _12138_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12069_ _09805_/A _12064_/X _09916_/A _12065_/X vssd1 vssd1 vccd1 vccd1 _12069_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_26_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06630_ _06627_/X _06629_/X _06627_/X _06629_/X vssd1 vssd1 vccd1 vccd1 _06630_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06561_ _06561_/A vssd1 vssd1 vccd1 vccd1 _06561_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08300_ _13922_/Q _08293_/X _08130_/X _08294_/X _08297_/X vssd1 vssd1 vccd1 vccd1
+ _13922_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09280_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09280_/X sky130_fd_sc_hd__clkbuf_2
X_06492_ _14639_/Q _09512_/A vssd1 vssd1 vccd1 vccd1 _06492_/Y sky130_fd_sc_hd__nand2_2
XFILLER_146_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ _08162_/A vssd1 vssd1 vccd1 vccd1 _08162_/X sky130_fd_sc_hd__buf_4
XFILLER_18_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07113_ _14510_/Q _07111_/X _06753_/X _07112_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _14510_/D sky130_fd_sc_hd__o221a_1
X_08093_ _08176_/A vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__inv_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07044_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ _08995_/A vssd1 vssd1 vccd1 vccd1 _08995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07946_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07877_ _14131_/Q _07808_/A _07876_/X _07811_/A _07872_/X vssd1 vssd1 vccd1 vccd1
+ _14131_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _09611_/X _09615_/X _09611_/X _09615_/X vssd1 vssd1 vccd1 vccd1 _09616_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06828_ _14606_/Q _06823_/X _06532_/X _08259_/A _06821_/X vssd1 vssd1 vccd1 vccd1
+ _14606_/D sky130_fd_sc_hd__o221a_1
XFILLER_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06759_ _08922_/A vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__buf_4
X_09547_ _09547_/A _12382_/X vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__and2_1
XFILLER_77_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _13277_/Q _09472_/X _12272_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _13277_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ _13851_/Q _08425_/X _08114_/X _08427_/X _08421_/X vssd1 vssd1 vccd1 vccd1
+ _13851_/D sky130_fd_sc_hd__o221a_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _14390_/Q vssd1 vssd1 vccd1 vccd1 _11440_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11371_ _13524_/Q vssd1 vssd1 vccd1 vccd1 _11371_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10322_ _14328_/Q vssd1 vssd1 vccd1 vccd1 _10322_/Y sky130_fd_sc_hd__inv_2
X_13110_ _13109_/X _12633_/X _13110_/S vssd1 vssd1 vccd1 vccd1 _13110_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14090_ _14169_/CLK _14090_/D vssd1 vssd1 vccd1 vccd1 _14090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13041_ _12600_/X _13040_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10253_ _10240_/Y _10242_/X _10243_/Y _10245_/X _10252_/X vssd1 vssd1 vccd1 vccd1
+ _10254_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10184_ _10184_/A vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13943_ _14100_/CLK _13943_/D vssd1 vssd1 vccd1 vccd1 _13943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13874_ _14107_/CLK _13874_/D vssd1 vssd1 vccd1 vccd1 _13874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12825_ _10048_/X _12824_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12825_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12756_ _09554_/X input338/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__mux2_1
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _14240_/Q _10696_/A _14435_/Q _10697_/A _11706_/X vssd1 vssd1 vccd1 vccd1
+ _11740_/B sky130_fd_sc_hd__a221oi_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12687_ _09591_/X _12686_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13194_/D sky130_fd_sc_hd__mux2_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14426_ _14595_/CLK _14426_/D vssd1 vssd1 vccd1 vccd1 _14426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11638_ _13647_/Q vssd1 vssd1 vccd1 vccd1 _11638_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14357_ _14629_/CLK _14357_/D vssd1 vssd1 vccd1 vccd1 _14357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ _13567_/Q _11430_/X _13808_/Q _11431_/X vssd1 vssd1 vccd1 vccd1 _11569_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13372_/CLK _13308_/D vssd1 vssd1 vccd1 vccd1 _13308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14288_ _14325_/CLK _14288_/D vssd1 vssd1 vccd1 vccd1 _14288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ _13368_/CLK _13239_/D vssd1 vssd1 vccd1 vccd1 _13271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07800_ _08190_/A vssd1 vssd1 vccd1 vccd1 _07800_/X sky130_fd_sc_hd__buf_4
X_08780_ _13677_/Q _08775_/X _08532_/X _08776_/X _08777_/X vssd1 vssd1 vccd1 vccd1
+ _13677_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07731_ _14199_/Q _07718_/X _07728_/X _07721_/X _07730_/X vssd1 vssd1 vccd1 vccd1
+ _14199_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07662_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07662_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09401_ _09401_/A _13091_/X vssd1 vssd1 vccd1 vccd1 _13333_/D sky130_fd_sc_hd__and2_1
X_06613_ _06614_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07593_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07593_/X sky130_fd_sc_hd__buf_2
XFILLER_129_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _13388_/Q _09326_/X _08181_/A _09327_/X _09330_/X vssd1 vssd1 vccd1 vccd1
+ _13388_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06544_ _06546_/A vssd1 vssd1 vccd1 vccd1 _06544_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _13427_/Q _09257_/X _08977_/X _09258_/X _09260_/X vssd1 vssd1 vccd1 vccd1
+ _13427_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08214_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08214_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09194_ _13466_/Q _09188_/X _08977_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1
+ _13466_/D sky130_fd_sc_hd__o221a_1
XFILLER_18_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08145_ _13995_/Q _08136_/X _08144_/X _08138_/X _08134_/X vssd1 vssd1 vccd1 vccd1
+ _13995_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08076_ _14024_/Q _08069_/X _07778_/X _08070_/X _08075_/X vssd1 vssd1 vccd1 vccd1
+ _14024_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07027_ _07062_/A vssd1 vssd1 vccd1 vccd1 _07027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput305 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _06493_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput316 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _06494_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput327 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _06503_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput338 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input338/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08978_ _13583_/Q _08969_/X _08977_/X _08971_/X _08975_/X vssd1 vssd1 vccd1 vccd1
+ _13583_/D sky130_fd_sc_hd__o221a_1
Xinput349 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 input349/X sky130_fd_sc_hd__buf_6
XFILLER_29_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07929_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10940_ _11412_/A vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__buf_2
XPHY_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10871_ _10869_/Y _10739_/X _10870_/Y _10741_/X vssd1 vssd1 vccd1 vccd1 _10871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12610_ _13324_/Q _12609_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13590_ _14188_/CLK _13590_/D vssd1 vssd1 vccd1 vccd1 _13590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12541_ _13375_/Q _10009_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__mux2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12472_ _12471_/X _06946_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__mux2_2
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14211_ _14325_/CLK _14211_/D vssd1 vssd1 vccd1 vccd1 _14211_/Q sky130_fd_sc_hd__dfxtp_1
X_11423_ _14000_/Q vssd1 vssd1 vccd1 vccd1 _11423_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_9 _11229_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _14183_/CLK _14142_/D vssd1 vssd1 vccd1 vccd1 _14142_/Q sky130_fd_sc_hd__dfxtp_1
X_11354_ _11354_/A _11354_/B _11354_/C _11354_/D vssd1 vssd1 vccd1 vccd1 _11354_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10305_ _11042_/A vssd1 vssd1 vccd1 vccd1 _10305_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14073_ _14459_/CLK _14073_/D vssd1 vssd1 vccd1 vccd1 _14073_/Q sky130_fd_sc_hd__dfxtp_1
X_11285_ _13841_/Q vssd1 vssd1 vccd1 vccd1 _11285_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10236_ _11685_/A vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _12592_/X input353/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13024_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10167_ _10697_/A vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10098_ _10098_/A _10132_/A vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__or2_1
XFILLER_97_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _14139_/CLK _13926_/D vssd1 vssd1 vccd1 vccd1 _13926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _14095_/CLK _13857_/D vssd1 vssd1 vccd1 vccd1 _13857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12808_ _12514_/X input356/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ _14121_/CLK _13788_/D vssd1 vssd1 vccd1 vccd1 _13788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12739_ _09541_/X _12738_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13213_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14409_ _14529_/CLK _14409_/D vssd1 vssd1 vccd1 vccd1 _14409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09950_ _09893_/A _09893_/B _09949_/Y vssd1 vssd1 vccd1 vccd1 _09950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08901_ _13614_/Q _08894_/X _08825_/X _08897_/X _08900_/X vssd1 vssd1 vccd1 vccd1
+ _13614_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _13287_/Q vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__inv_2
XFILLER_154_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08832_ _08868_/A vssd1 vssd1 vccd1 vccd1 _08832_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08763_ _13688_/Q _08758_/X _08505_/X _08760_/X _08761_/X vssd1 vssd1 vccd1 vccd1
+ _13688_/D sky130_fd_sc_hd__o221a_1
XPHY_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07714_ _07714_/A vssd1 vssd1 vccd1 vccd1 _07714_/X sky130_fd_sc_hd__buf_4
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__buf_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07645_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__buf_4
XPHY_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07576_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07576_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06527_ _08660_/A _11673_/A vssd1 vssd1 vccd1 vccd1 _06811_/A sky130_fd_sc_hd__or2_2
XFILLER_107_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _13399_/Q _09310_/X _08155_/A _09311_/X _09314_/X vssd1 vssd1 vccd1 vccd1
+ _13399_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09246_ _13438_/Q _09241_/X _08950_/X _09242_/X _09244_/X vssd1 vssd1 vccd1 vccd1
+ _13438_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ _13476_/Q _09171_/X _09035_/X _09172_/X _09173_/X vssd1 vssd1 vccd1 vccd1
+ _13476_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08128_ _08128_/A vssd1 vssd1 vccd1 vccd1 _08128_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08059_ _14034_/Q _08053_/X _07753_/X _08054_/X _08058_/X vssd1 vssd1 vccd1 vccd1
+ _14034_/D sky130_fd_sc_hd__o221a_1
XFILLER_150_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11070_ _13914_/Q vssd1 vssd1 vccd1 vccd1 _11070_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10021_ _13379_/Q _10020_/B _10022_/A vssd1 vssd1 vccd1 vccd1 _10021_/X sky130_fd_sc_hd__o21a_1
Xinput102 la_data_in[41] vssd1 vssd1 vccd1 vccd1 _06603_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput113 la_data_in[51] vssd1 vssd1 vccd1 vccd1 _06668_/A sky130_fd_sc_hd__buf_2
XPHY_7134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput124 la_data_in[61] vssd1 vssd1 vccd1 vccd1 _06545_/A sky130_fd_sc_hd__buf_2
XFILLER_27_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput135 la_data_in[71] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__buf_1
XPHY_7156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 la_data_in[81] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__buf_1
XPHY_7167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 la_data_in[91] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__buf_1
XPHY_7178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 la_oenb[100] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__buf_1
XPHY_7189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 la_oenb[110] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__buf_1
XFILLER_40_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _14636_/Q vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__inv_2
XPHY_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _14146_/CLK _13711_/D vssd1 vssd1 vccd1 vccd1 _13711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10923_ _11397_/A vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13642_ _14143_/CLK _13642_/D vssd1 vssd1 vccd1 vccd1 _13642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10854_ _10852_/Y _10709_/X _10853_/Y _10711_/X vssd1 vssd1 vccd1 vccd1 _10854_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13573_ _14130_/CLK _13573_/D vssd1 vssd1 vccd1 vccd1 _13573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10785_ _13589_/Q vssd1 vssd1 vccd1 vccd1 _10785_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _13360_/Q _10039_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12524_/X sky130_fd_sc_hd__mux2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12455_ _12509_/X _06927_/Y _12455_/S vssd1 vssd1 vccd1 vccd1 _12455_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11406_ _11406_/A vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__clkbuf_4
X_12386_ _13209_/Q _08945_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__mux2_1
X_14125_ _14130_/CLK _14125_/D vssd1 vssd1 vccd1 vccd1 _14125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11337_ _14622_/Q vssd1 vssd1 vccd1 vccd1 _11337_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _14056_/CLK _14056_/D vssd1 vssd1 vccd1 vccd1 _14056_/Q sky130_fd_sc_hd__dfxtp_1
X_11268_ _11266_/Y _11223_/X _11267_/Y _11225_/X vssd1 vssd1 vccd1 vccd1 _11268_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13007_ _12582_/X _13006_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__mux2_1
X_10219_ _11673_/A vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _14143_/CLK _13909_/D vssd1 vssd1 vccd1 vccd1 _13909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07430_ _14356_/Q _07422_/X _07330_/X _07424_/X _07425_/X vssd1 vssd1 vccd1 vccd1
+ _14356_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07361_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07361_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _13520_/Q _09095_/X _08940_/X _09096_/X _09093_/X vssd1 vssd1 vccd1 vccd1
+ _13520_/D sky130_fd_sc_hd__o221a_1
X_07292_ _14412_/Q _07290_/X _06825_/X _07291_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _14412_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09933_ _13304_/Q _09931_/Y _09899_/B vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09864_ _13304_/Q vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__inv_2
XFILLER_86_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08815_ _09132_/A _11639_/A vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__or2_2
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09793_/A _09793_/B _09794_/Y vssd1 vssd1 vccd1 vccd1 _09795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _08801_/A vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__inv_2
XPHY_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_207 _13275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08677_/A vssd1 vssd1 vccd1 vccd1 _08677_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07628_ _08989_/A vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ _07614_/A vssd1 vssd1 vccd1 vccd1 _07613_/A sky130_fd_sc_hd__inv_2
XFILLER_165_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ _14216_/Q _10437_/X _14411_/Q _10438_/X _10569_/X vssd1 vssd1 vccd1 vccd1
+ _10603_/B sky130_fd_sc_hd__a221oi_2
XFILLER_210_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09229_ _13449_/Q _09224_/X _08920_/X _09225_/X _09228_/X vssd1 vssd1 vccd1 vccd1
+ _13449_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12240_ _12240_/A vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12171_ vssd1 vssd1 vccd1 vccd1 _12171_/HI _12171_/LO sky130_fd_sc_hd__conb_1
XFILLER_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11122_ _13636_/Q vssd1 vssd1 vccd1 vccd1 _11122_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11053_ _13517_/Q vssd1 vssd1 vccd1 vccd1 _11053_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10004_ _13373_/Q _10004_/B vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _14246_/Q _11830_/X _14441_/Q _11831_/X vssd1 vssd1 vccd1 vccd1 _11955_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10906_ _10904_/Y _10729_/X _10905_/Y _10731_/X vssd1 vssd1 vccd1 vccd1 _10906_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11886_ _13574_/Q _10206_/A _13815_/Q _10209_/A vssd1 vssd1 vccd1 vccd1 _11886_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13625_ _14047_/CLK _13625_/D vssd1 vssd1 vccd1 vccd1 _13625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10837_ _10832_/Y _10745_/X _10833_/Y _10747_/X _10836_/X vssd1 vssd1 vccd1 vccd1
+ _10838_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13556_ _14114_/CLK _13556_/D vssd1 vssd1 vccd1 vccd1 _13556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ _13830_/Q vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12507_ _12506_/X _10057_/Y _12507_/S vssd1 vssd1 vccd1 vccd1 _12507_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13487_ _14470_/CLK _13487_/D vssd1 vssd1 vccd1 vccd1 _13487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10699_ _13393_/Q _10568_/X _13705_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _10699_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _12437_/X _06906_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12438_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput406 _12076_/LO vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput417 _12077_/LO vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput428 _12078_/LO vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput439 _12081_/LO vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12369_ _13199_/Q _12368_/X input78/X vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14108_ _14110_/CLK _14108_/D vssd1 vssd1 vccd1 vccd1 _14108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14039_ _14119_/CLK _14039_/D vssd1 vssd1 vccd1 vccd1 _14039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06930_ _14580_/Q vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06861_ _06861_/A vssd1 vssd1 vccd1 vccd1 _06861_/X sky130_fd_sc_hd__buf_1
XFILLER_110_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08600_ _08644_/A vssd1 vssd1 vccd1 vccd1 _08636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09580_ _09586_/A _12325_/X vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__and2_1
X_06792_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08531_ _13802_/Q _08526_/X _08530_/X _08528_/X _08524_/X vssd1 vssd1 vccd1 vccd1
+ _13802_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08462_ _13832_/Q _08460_/X _08162_/X _08461_/X _08457_/X vssd1 vssd1 vccd1 vccd1
+ _13832_/D sky130_fd_sc_hd__o221a_1
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07413_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__clkbuf_2
X_08393_ _13869_/Q _08388_/X _08167_/X _08389_/X _08392_/X vssd1 vssd1 vccd1 vccd1
+ _13869_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07344_ _14390_/Q _07335_/X _07343_/X _07337_/X _07333_/X vssd1 vssd1 vccd1 vccd1
+ _14390_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07275_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07275_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09039_/A vssd1 vssd1 vccd1 vccd1 _09014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__or2_2
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _13080_/S sky130_fd_sc_hd__and2_4
XFILLER_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09778_ _09778_/A _09833_/A vssd1 vssd1 vccd1 vccd1 _09779_/B sky130_fd_sc_hd__or2_1
XFILLER_74_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _13704_/Q _08722_/X _08562_/X _08723_/X _08728_/X vssd1 vssd1 vccd1 vccd1
+ _13704_/D sky130_fd_sc_hd__o221a_1
XPHY_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11740_ _11740_/A _11740_/B _11740_/C _11740_/D vssd1 vssd1 vccd1 vccd1 _11740_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A vssd1 vssd1 vccd1 vccd1 _11671_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13410_ _14183_/CLK _13410_/D vssd1 vssd1 vccd1 vccd1 _13410_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10622_ _10612_/Y _10445_/X _10615_/X _10618_/X _10621_/X vssd1 vssd1 vccd1 vccd1
+ _10644_/C sky130_fd_sc_hd__o2111a_4
X_14390_ _14629_/CLK _14390_/D vssd1 vssd1 vccd1 vccd1 _14390_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13341_ _14538_/CLK _13341_/D vssd1 vssd1 vccd1 vccd1 _13341_/Q sky130_fd_sc_hd__dfxtp_1
X_10553_ _10548_/Y _10492_/X _10549_/Y _10495_/X _10552_/X vssd1 vssd1 vccd1 vccd1
+ _10560_/C sky130_fd_sc_hd__o221a_1
XFILLER_13_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13272_ _13368_/CLK _13272_/D vssd1 vssd1 vccd1 vccd1 _13272_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10484_ _11439_/A vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12154_ vssd1 vssd1 vccd1 vccd1 _12154_/HI _12154_/LO sky130_fd_sc_hd__conb_1
XFILLER_174_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ _14305_/Q vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12085_ vssd1 vssd1 vccd1 vccd1 _12085_/HI _12085_/LO sky130_fd_sc_hd__conb_1
XFILLER_81_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11036_ _14070_/Q vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ _12572_/X _12986_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12987_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11938_ _14284_/Q vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11869_ _13691_/Q vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13608_ _14481_/CLK _13608_/D vssd1 vssd1 vccd1 vccd1 _13608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14588_ _14621_/CLK _14588_/D vssd1 vssd1 vccd1 vccd1 _14588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13539_ _14123_/CLK _13539_/D vssd1 vssd1 vccd1 vccd1 _13539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07060_ _14535_/Q _07052_/X _06801_/X _07053_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _14535_/D sky130_fd_sc_hd__o221a_1
XFILLER_199_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07962_ _14088_/Q _07955_/X _07712_/X _07957_/X _07960_/X vssd1 vssd1 vccd1 vccd1
+ _14088_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _09701_/A vssd1 vssd1 vccd1 vccd1 _09701_/Y sky130_fd_sc_hd__inv_2
X_06913_ _06901_/X _12297_/X _06912_/Y _06903_/X vssd1 vssd1 vccd1 vccd1 _06914_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_190_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07893_ _07935_/A vssd1 vssd1 vccd1 vccd1 _07927_/A sky130_fd_sc_hd__buf_4
XFILLER_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09632_ _06889_/Y _14581_/Q _14591_/Q _06927_/Y vssd1 vssd1 vccd1 vccd1 _09632_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06844_ _08983_/A vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ _09573_/A _12352_/X vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__and2_1
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06775_ _08140_/A vssd1 vssd1 vccd1 vccd1 _06775_/X sky130_fd_sc_hd__buf_2
XFILLER_208_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _08917_/A vssd1 vssd1 vccd1 vccd1 _08514_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09494_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _13879_/Q _08371_/X _08142_/X _08372_/X _08375_/X vssd1 vssd1 vccd1 vccd1
+ _13879_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07327_ _07723_/A vssd1 vssd1 vccd1 vccd1 _07327_/X sky130_fd_sc_hd__buf_2
XFILLER_143_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07189_ _07213_/A vssd1 vssd1 vccd1 vccd1 _07189_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12910_ _12538_/X _12909_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13890_ _14100_/CLK _13890_/D vssd1 vssd1 vccd1 vccd1 _13890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12841_ _12521_/X _12840_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12772_ _09522_/X input351/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__mux2_1
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14511_ _14629_/CLK _14511_/D vssd1 vssd1 vccd1 vccd1 _14511_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11723_ _14630_/Q vssd1 vssd1 vccd1 vccd1 _11723_/Y sky130_fd_sc_hd__inv_2
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14442_ _14481_/CLK _14442_/D vssd1 vssd1 vccd1 vccd1 _14442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11654_ _14122_/Q vssd1 vssd1 vccd1 vccd1 _11654_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10605_ _13430_/Q vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__inv_2
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14373_ _14629_/CLK _14373_/D vssd1 vssd1 vccd1 vccd1 _14373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11585_ _13489_/Q vssd1 vssd1 vccd1 vccd1 _11585_/Y sky130_fd_sc_hd__inv_2
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13324_ _13877_/CLK _13324_/D vssd1 vssd1 vccd1 vccd1 _13324_/Q sky130_fd_sc_hd__dfxtp_1
X_10536_ _13506_/Q vssd1 vssd1 vccd1 vccd1 _10536_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13255_ _13352_/CLK _13255_/D vssd1 vssd1 vccd1 vccd1 _13255_/Q sky130_fd_sc_hd__dfxtp_4
X_10467_ _10443_/Y _10445_/X _10452_/X _10459_/X _10466_/X vssd1 vssd1 vccd1 vccd1
+ _10519_/C sky130_fd_sc_hd__o2111a_4
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13186_ _14573_/Q _14574_/Q _14571_/Q _14572_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13186_/X sky130_fd_sc_hd__mux4_1
X_10398_ _13504_/Q vssd1 vssd1 vccd1 vccd1 _10398_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12137_ vssd1 vssd1 vccd1 vccd1 _12137_/HI _12137_/LO sky130_fd_sc_hd__conb_1
XFILLER_65_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12068_ _09801_/A _12064_/X _09912_/A _12065_/X vssd1 vssd1 vccd1 vccd1 _12068_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_93_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _14381_/Q vssd1 vssd1 vccd1 vccd1 _11019_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06560_ _06556_/Y _08960_/A _08954_/A _06559_/Y vssd1 vssd1 vccd1 vccd1 _06561_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_59_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06491_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06918_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_146_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08230_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07112_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08092_ _08341_/A _11658_/A vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__or2_4
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07043_ _14545_/Q _07035_/X _06766_/X _07036_/X _07038_/X vssd1 vssd1 vccd1 vccd1
+ _14545_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ _09049_/A vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07945_ _14095_/Q _07882_/A _07796_/X _07884_/A _07940_/X vssd1 vssd1 vccd1 vccd1
+ _14095_/D sky130_fd_sc_hd__o221a_1
XPHY_6818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07876_ _08268_/A vssd1 vssd1 vccd1 vccd1 _07876_/X sky130_fd_sc_hd__buf_4
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _09612_/X _09614_/X _09612_/X _09614_/X vssd1 vssd1 vccd1 vccd1 _09615_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06827_ _09051_/A vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__buf_4
X_09546_ _09544_/X _09543_/X _13276_/Q _09545_/X vssd1 vssd1 vccd1 vccd1 _13244_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06758_ _14626_/Q _06751_/X _06757_/X _06754_/X _06749_/X vssd1 vssd1 vccd1 vccd1
+ _14626_/D sky130_fd_sc_hd__o221a_1
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _13278_/Q _09472_/X _12273_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _13278_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _06682_/Y _06688_/X _06682_/Y _06688_/X vssd1 vssd1 vccd1 vccd1 _06691_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_184_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ _13852_/Q _08425_/X _08110_/X _08427_/X _08421_/X vssd1 vssd1 vccd1 vccd1
+ _13852_/D sky130_fd_sc_hd__o221a_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08359_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08359_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _13999_/Q vssd1 vssd1 vccd1 vccd1 _11370_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _14484_/Q vssd1 vssd1 vccd1 vccd1 _10321_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13040_ _12600_/X input348/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13040_/X sky130_fd_sc_hd__mux2_1
X_10252_ _10246_/Y _10248_/X _10249_/Y _10251_/X vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10183_ _11650_/A vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13942_ _14100_/CLK _13942_/D vssd1 vssd1 vccd1 vccd1 _13942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13873_ _14107_/CLK _13873_/D vssd1 vssd1 vccd1 vccd1 _13873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12824_ _10048_/X input330/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12755_ _09552_/X _12754_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13209_/D sky130_fd_sc_hd__mux2_1
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _13414_/Q _11514_/X _13726_/Q _11642_/X vssd1 vssd1 vccd1 vccd1 _11706_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12686_ _09591_/X _12685_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12686_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14621_/CLK _14425_/D vssd1 vssd1 vccd1 vccd1 _14425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__buf_2
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14629_/CLK _14356_/D vssd1 vssd1 vccd1 vccd1 _14356_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11568_ _11558_/Y _11412_/X _11561_/X _11564_/X _11567_/X vssd1 vssd1 vccd1 vccd1
+ _11590_/C sky130_fd_sc_hd__o2111a_4
XFILLER_144_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13307_ _13371_/CLK _13307_/D vssd1 vssd1 vccd1 vccd1 _13307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10519_ _10519_/A _10519_/B _10519_/C _10519_/D vssd1 vssd1 vccd1 vccd1 _10519_/Y
+ sky130_fd_sc_hd__nand4_4
X_14287_ _14325_/CLK _14287_/D vssd1 vssd1 vccd1 vccd1 _14287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11499_ _11494_/Y _11445_/X _11495_/Y _11447_/X _11498_/X vssd1 vssd1 vccd1 vccd1
+ _11506_/C sky130_fd_sc_hd__o221a_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13238_ _13368_/CLK _13238_/D vssd1 vssd1 vccd1 vccd1 _13270_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13169_ _12663_/X _13168_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07730_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07730_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07661_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07661_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09400_ _09401_/A _13087_/X vssd1 vssd1 vccd1 vccd1 _13334_/D sky130_fd_sc_hd__and2_1
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06612_ _06573_/X _06561_/A _08912_/A _06561_/Y vssd1 vssd1 vccd1 vccd1 _06612_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07592_ _14270_/Q _07589_/X _07352_/X _07590_/X _07585_/X vssd1 vssd1 vccd1 vccd1
+ _14270_/D sky130_fd_sc_hd__o221a_1
XFILLER_207_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _13389_/Q _09326_/X _08179_/A _09327_/X _09330_/X vssd1 vssd1 vccd1 vccd1
+ _13389_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06543_ _06545_/A vssd1 vssd1 vccd1 vccd1 _08827_/A sky130_fd_sc_hd__buf_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09262_ _13428_/Q _09257_/X _08974_/X _09258_/X _09260_/X vssd1 vssd1 vccd1 vccd1
+ _13428_/D sky130_fd_sc_hd__o221a_1
XFILLER_90_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08213_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08213_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09193_ _13467_/Q _09188_/X _08974_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1
+ _13467_/D sky130_fd_sc_hd__o221a_1
XFILLER_72_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08144_ _08144_/A vssd1 vssd1 vccd1 vccd1 _08144_/X sky130_fd_sc_hd__buf_4
XFILLER_159_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08075_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07026_ _07070_/A vssd1 vssd1 vccd1 vccd1 _07062_/A sky130_fd_sc_hd__buf_4
XFILLER_66_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput306 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _06493_/D sky130_fd_sc_hd__clkbuf_1
XPHY_7327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput317 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input317/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08977_ _08977_/A vssd1 vssd1 vccd1 vccd1 _08977_/X sky130_fd_sc_hd__buf_4
Xinput328 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _06503_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput339 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input339/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07928_ _14105_/Q _07926_/X _07771_/X _07927_/X _07921_/X vssd1 vssd1 vccd1 vccd1
+ _14105_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07859_ _14143_/Q _07855_/X _07774_/X _07856_/X _07857_/X vssd1 vssd1 vccd1 vccd1
+ _14143_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10870_ _14261_/Q vssd1 vssd1 vccd1 vccd1 _10870_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09583_/A vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _13376_/Q _10012_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12540_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12471_ _12470_/X _06946_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12471_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ _14325_/CLK _14210_/D vssd1 vssd1 vccd1 vccd1 _14210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11422_ _11418_/Y _11419_/X _11420_/Y _11421_/X vssd1 vssd1 vccd1 vccd1 _11422_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14141_ _14143_/CLK _14141_/D vssd1 vssd1 vccd1 vccd1 _14141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11353_ _11334_/X _11353_/B _11353_/C _11353_/D vssd1 vssd1 vccd1 vccd1 _11354_/D
+ sky130_fd_sc_hd__and4b_1
X_10304_ _10299_/Y _10150_/X _10300_/Y _10153_/X _10303_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/A sky130_fd_sc_hd__o221a_2
XFILLER_141_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14072_ _14188_/CLK _14072_/D vssd1 vssd1 vccd1 vccd1 _14072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ _11282_/Y _11178_/X _11283_/Y _11180_/X vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13023_ _12590_/X _13022_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13023_/X sky130_fd_sc_hd__mux2_1
X_10235_ _14248_/Q vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10166_ _11831_/A vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10097_ _10097_/A _12478_/X vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__nor2_8
XFILLER_43_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13925_ _14119_/CLK _13925_/D vssd1 vssd1 vccd1 vccd1 _13925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13856_ _14095_/CLK _13856_/D vssd1 vssd1 vccd1 vccd1 _13856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _12513_/X _12806_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12807_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13787_ _14121_/CLK _13787_/D vssd1 vssd1 vccd1 vccd1 _13787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ _10994_/Y _10923_/X _10995_/Y _10925_/X _10998_/X vssd1 vssd1 vccd1 vccd1
+ _11035_/A sky130_fd_sc_hd__o221a_2
XFILLER_128_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12738_ _09541_/X _12737_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12738_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _09580_/X _12668_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12669_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ _14481_/CLK _14408_/D vssd1 vssd1 vccd1 vccd1 _14408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14339_ _14611_/CLK _14339_/D vssd1 vssd1 vccd1 vccd1 _14339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08900_ _08923_/A vssd1 vssd1 vccd1 vccd1 _08900_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09880_ _13288_/Q vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__inv_2
XFILLER_48_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08831_ _08876_/A vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08762_ _13689_/Q _08758_/X _08501_/X _08760_/X _08761_/X vssd1 vssd1 vccd1 vccd1
+ _13689_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07713_ _14205_/Q _07704_/X _07712_/X _07706_/X _07698_/X vssd1 vssd1 vccd1 vccd1
+ _14205_/D sky130_fd_sc_hd__o221a_1
X_08693_ _13725_/Q _08687_/X _08508_/X _08689_/X _08684_/X vssd1 vssd1 vccd1 vccd1
+ _13725_/D sky130_fd_sc_hd__o221a_1
XPHY_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07644_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07575_ _14280_/Q _07571_/X _07327_/X _07573_/X _07566_/X vssd1 vssd1 vccd1 vccd1
+ _14280_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09314_ _09519_/A vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__clkbuf_2
X_06526_ _07803_/A _09271_/B _08989_/C _09271_/D vssd1 vssd1 vccd1 vccd1 _11673_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_107_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _13439_/Q _09241_/X _08948_/X _09242_/X _09244_/X vssd1 vssd1 vccd1 vccd1
+ _13439_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _13477_/Q _09171_/X _08950_/X _09172_/X _09173_/X vssd1 vssd1 vccd1 vccd1
+ _13477_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08127_ _14002_/Q _08122_/X _08126_/X _08124_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _14002_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08058_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07009_ _08989_/D vssd1 vssd1 vccd1 vccd1 _07630_/D sky130_fd_sc_hd__buf_1
XFILLER_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10020_ _13379_/Q _10020_/B vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput103 la_data_in[42] vssd1 vssd1 vccd1 vccd1 _06558_/A sky130_fd_sc_hd__buf_2
XFILLER_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput114 la_data_in[52] vssd1 vssd1 vccd1 vccd1 _06565_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 la_data_in[62] vssd1 vssd1 vccd1 vccd1 _06541_/A sky130_fd_sc_hd__buf_2
XPHY_7146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 la_data_in[72] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__buf_1
XPHY_7157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput147 la_data_in[82] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__buf_1
XPHY_7168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 la_data_in[92] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__buf_1
XPHY_7179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 la_oenb[101] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__buf_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _14363_/Q vssd1 vssd1 vccd1 vccd1 _11971_/Y sky130_fd_sc_hd__inv_2
XPHY_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13710_ _14146_/CLK _13710_/D vssd1 vssd1 vccd1 vccd1 _13710_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10922_ _14068_/Q vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__inv_2
XPHY_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13641_ _14143_/CLK _13641_/D vssd1 vssd1 vccd1 vccd1 _13641_/Q sky130_fd_sc_hd__dfxtp_1
X_10853_ _14105_/Q vssd1 vssd1 vccd1 vccd1 _10853_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _14123_/CLK _13572_/D vssd1 vssd1 vccd1 vccd1 _13572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10784_ _14298_/Q vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _13361_/Q _10040_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12454_ _12453_/X _06924_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11405_ _11396_/Y _11397_/X _11398_/Y _11399_/X _11404_/X vssd1 vssd1 vccd1 vccd1
+ _11465_/A sky130_fd_sc_hd__o221a_2
XFILLER_201_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12385_ _12384_/X _13210_/Q _12645_/S vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__mux2_1
X_14124_ _14130_/CLK _14124_/D vssd1 vssd1 vccd1 vccd1 _14124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11336_ _14349_/Q vssd1 vssd1 vccd1 vccd1 _11336_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14055_ _14056_/CLK _14055_/D vssd1 vssd1 vccd1 vccd1 _14055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11267_ _14464_/Q vssd1 vssd1 vccd1 vccd1 _11267_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13006_ _13005_/X _12582_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10218_ _14599_/Q vssd1 vssd1 vccd1 vccd1 _10218_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11198_ _14502_/Q vssd1 vssd1 vccd1 vccd1 _11198_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _11633_/A vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _14143_/CLK _13908_/D vssd1 vssd1 vccd1 vccd1 _13908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13839_ _13996_/CLK _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07360_ _14384_/Q _07348_/X _07358_/X _07350_/X _07359_/X vssd1 vssd1 vccd1 vccd1
+ _14384_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ _09039_/A vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ _09897_/A _09897_/B _09931_/Y vssd1 vssd1 vccd1 vccd1 _09932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09863_ _13305_/Q vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__inv_2
XFILLER_8_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08814_ _08814_/A _08890_/B _08814_/C _09201_/D vssd1 vssd1 vccd1 vccd1 _11639_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_41_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09794_ _09798_/B vssd1 vssd1 vccd1 vccd1 _09794_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08745_ _08745_/A _11637_/A vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__or2_2
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _13276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08676_ _08730_/A vssd1 vssd1 vccd1 vccd1 _08677_/A sky130_fd_sc_hd__buf_2
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07627_ _09272_/A vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__buf_4
XPHY_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _07558_/A _11685_/A vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__or2_2
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ _09458_/A _09511_/A _06509_/C vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__or3_4
XFILLER_194_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07489_ _07542_/A vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09228_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__buf_2
XFILLER_127_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _13488_/Q _09155_/X _08920_/X _09156_/X _09157_/X vssd1 vssd1 vccd1 vccd1
+ _13488_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12170_ vssd1 vssd1 vccd1 vccd1 _12170_/HI _12170_/LO sky130_fd_sc_hd__conb_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _13675_/Q vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11052_ _13992_/Q vssd1 vssd1 vccd1 vccd1 _11052_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _10003_/A vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__inv_2
XFILLER_153_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11954_ _11949_/Y _10150_/A _11950_/Y _10153_/A _11953_/X vssd1 vssd1 vccd1 vccd1
+ _11989_/A sky130_fd_sc_hd__o221a_2
XPHY_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _14379_/Q vssd1 vssd1 vccd1 vccd1 _10905_/Y sky130_fd_sc_hd__inv_2
XPHY_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11885_ _11875_/Y _10178_/A _11878_/X _11881_/X _11884_/X vssd1 vssd1 vccd1 vccd1
+ _11907_/C sky130_fd_sc_hd__o2111a_4
XPHY_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13624_ _14047_/CLK _13624_/D vssd1 vssd1 vccd1 vccd1 _13624_/Q sky130_fd_sc_hd__dfxtp_1
X_10836_ _10834_/Y _10749_/X _10835_/Y _10751_/X vssd1 vssd1 vccd1 vccd1 _10836_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _14114_/CLK _13555_/D vssd1 vssd1 vccd1 vccd1 _13555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10767_ _10765_/Y _10704_/X _10766_/Y _10706_/X vssd1 vssd1 vccd1 vccd1 _10767_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12506_ _14561_/Q _14562_/Q _12506_/S vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13486_ _14470_/CLK _13486_/D vssd1 vssd1 vccd1 vccd1 _13486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10698_ _11408_/A vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12509_/X _06906_/Y _12437_/S vssd1 vssd1 vccd1 vccd1 _12437_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput407 _12086_/LO vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput418 _12234_/A vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12368_ _13199_/Q input96/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__mux2_1
Xoutput429 _12244_/A vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14107_ _14107_/CLK _14107_/D vssd1 vssd1 vccd1 vccd1 _14107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11319_ _11314_/Y _11161_/X _11315_/Y _11163_/X _11318_/X vssd1 vssd1 vccd1 vccd1
+ _11354_/A sky130_fd_sc_hd__o221a_2
XFILLER_180_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12299_ _11354_/Y _14544_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14038_ _14119_/CLK _14038_/D vssd1 vssd1 vccd1 vccd1 _14038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06860_ _06976_/A vssd1 vssd1 vccd1 vccd1 _06861_/A sky130_fd_sc_hd__buf_1
XFILLER_110_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06791_ _14617_/Q _06787_/X _06789_/X _06790_/X _06785_/X vssd1 vssd1 vccd1 vccd1
+ _14617_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08530_ _08933_/A vssd1 vssd1 vccd1 vccd1 _08530_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_208_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08461_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08461_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07412_ _07809_/A vssd1 vssd1 vccd1 vccd1 _07412_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08392_ _08421_/A vssd1 vssd1 vccd1 vccd1 _08392_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07343_ _08130_/A vssd1 vssd1 vccd1 vccd1 _07343_/X sky130_fd_sc_hd__buf_2
XFILLER_36_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07274_ _07282_/A vssd1 vssd1 vccd1 vccd1 _07274_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09013_ _13568_/Q _09004_/X _08914_/X _09006_/X _09011_/X vssd1 vssd1 vccd1 vccd1
+ _13568_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _13371_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_172_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09915_ _13314_/Q vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__inv_2
XFILLER_99_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09846_ _13319_/Q _12634_/S _09770_/B _12233_/A vssd1 vssd1 vccd1 vccd1 _09846_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__or2_1
XFILLER_210_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06989_ _06989_/A vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08728_ _08728_/A vssd1 vssd1 vccd1 vccd1 _08728_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08659_ _09131_/A _09271_/B _09063_/C _08673_/D vssd1 vssd1 vccd1 vccd1 _09599_/A
+ sky130_fd_sc_hd__or4_4
XPHY_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11670_ _14356_/Q vssd1 vssd1 vccd1 vccd1 _11670_/Y sky130_fd_sc_hd__inv_2
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10619_/Y _10462_/X _10620_/Y _10465_/X vssd1 vssd1 vccd1 vccd1 _10621_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13340_ _13372_/CLK _13340_/D vssd1 vssd1 vccd1 vccd1 _13340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ _10550_/Y _10498_/X _10551_/Y _10501_/X vssd1 vssd1 vccd1 vccd1 _10552_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _13877_/CLK _13271_/D vssd1 vssd1 vccd1 vccd1 _13271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10483_ _11673_/A vssd1 vssd1 vccd1 vccd1 _11439_/A sky130_fd_sc_hd__buf_2
XFILLER_87_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12153_ vssd1 vssd1 vccd1 vccd1 _12153_/HI _12153_/LO sky130_fd_sc_hd__conb_1
XFILLER_151_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11104_ _11099_/Y _10963_/X _11100_/Y _10965_/X _11103_/X vssd1 vssd1 vccd1 vccd1
+ _11117_/B sky130_fd_sc_hd__o221a_2
XFILLER_46_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12084_ vssd1 vssd1 vccd1 vccd1 _12084_/HI _12084_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ _11035_/A _11035_/B _11035_/C _11035_/D vssd1 vssd1 vccd1 vccd1 _11035_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_42_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _12985_/X _12572_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11937_ _14206_/Q vssd1 vssd1 vccd1 vccd1 _11937_/Y sky130_fd_sc_hd__inv_2
XPHY_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11868_ _13457_/Q vssd1 vssd1 vccd1 vccd1 _11868_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _14481_/CLK _13607_/D vssd1 vssd1 vccd1 vccd1 _13607_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ _13203_/Q _10775_/X _14026_/Q _10719_/X _10818_/X vssd1 vssd1 vccd1 vccd1
+ _10819_/X sky130_fd_sc_hd__a221o_4
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ _13533_/Q vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14587_ _14621_/CLK _14587_/D vssd1 vssd1 vccd1 vccd1 _14587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13538_ _14130_/CLK _13538_/D vssd1 vssd1 vccd1 vccd1 _13538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13469_ _14178_/CLK _13469_/D vssd1 vssd1 vccd1 vccd1 _13469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ _14089_/Q _07955_/X _07710_/X _07957_/X _07960_/X vssd1 vssd1 vccd1 vccd1
+ _14089_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09700_ _06897_/X _14585_/Q _14589_/Q _06912_/Y vssd1 vssd1 vccd1 vccd1 _09701_/A
+ sky130_fd_sc_hd__o22a_1
X_06912_ _14585_/Q vssd1 vssd1 vccd1 vccd1 _06912_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07892_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09631_ _09629_/X _09630_/X _09629_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _09631_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06843_ _12396_/S _06843_/B vssd1 vssd1 vccd1 vccd1 _06843_/X sky130_fd_sc_hd__and2_1
XFILLER_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09562_ _09588_/A vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06774_ _08933_/A vssd1 vssd1 vccd1 vccd1 _08140_/A sky130_fd_sc_hd__buf_4
XFILLER_77_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08513_ _08552_/A vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09493_ _09500_/A vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _08460_/A vssd1 vssd1 vccd1 vccd1 _08444_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07326_ _14398_/Q _07322_/X _07323_/X _07325_/X _07319_/X vssd1 vssd1 vccd1 vccd1
+ _14398_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07257_ _07282_/A vssd1 vssd1 vccd1 vccd1 _07257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07188_ _14470_/Q _07185_/X _06757_/X _07186_/X _07181_/X vssd1 vssd1 vccd1 vccd1
+ _14470_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09829_ _13340_/Q _09827_/Y _09791_/B vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12840_ _12521_/X input333/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12771_ _09519_/X _12770_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13221_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _14357_/Q vssd1 vssd1 vccd1 vccd1 _11722_/Y sky130_fd_sc_hd__inv_2
X_14510_ _14629_/CLK _14510_/D vssd1 vssd1 vccd1 vccd1 _14510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _14481_/CLK _14441_/D vssd1 vssd1 vccd1 vccd1 _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _11653_/A vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10604_ _14061_/Q vssd1 vssd1 vccd1 vccd1 _10604_/Y sky130_fd_sc_hd__inv_2
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14372_ _14629_/CLK _14372_/D vssd1 vssd1 vccd1 vccd1 _14372_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11584_ _14159_/Q vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13323_ _13877_/CLK _13323_/D vssd1 vssd1 vccd1 vccd1 _13323_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ _13981_/Q vssd1 vssd1 vccd1 vccd1 _10535_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13254_ _13372_/CLK _13254_/D vssd1 vssd1 vccd1 vccd1 _13286_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10466_ _10460_/Y _10462_/X _10463_/Y _10465_/X vssd1 vssd1 vccd1 vccd1 _10466_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_178_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _14565_/Q _14566_/Q _14563_/Q _14564_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13185_/X sky130_fd_sc_hd__mux4_2
X_10397_ _13979_/Q vssd1 vssd1 vccd1 vccd1 _10397_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ vssd1 vssd1 vccd1 vccd1 _12136_/HI _12136_/LO sky130_fd_sc_hd__conb_1
XFILLER_170_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12067_ _09798_/A _12064_/X _09909_/A _12065_/X vssd1 vssd1 vccd1 vccd1 _12067_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_152_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ _14615_/Q vssd1 vssd1 vccd1 vccd1 _11018_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12564_/X _12968_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _12969_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06490_ _12282_/X vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _14639_/CLK _14639_/D vssd1 vssd1 vccd1 vccd1 _14639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08160_ _13989_/Q _08149_/X _08158_/X _08151_/X _08159_/X vssd1 vssd1 vccd1 vccd1
+ _13989_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07111_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _08411_/A _08890_/B _09271_/C _08091_/D vssd1 vssd1 vccd1 vccd1 _11658_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_200_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07042_ _14546_/Q _07035_/X _06763_/X _07036_/X _07038_/X vssd1 vssd1 vccd1 vccd1
+ _14546_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08993_ _08993_/A vssd1 vssd1 vccd1 vccd1 _08993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07944_ _14096_/Q _07934_/X _07792_/X _07935_/X _07940_/X vssd1 vssd1 vccd1 vccd1
+ _14096_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _14132_/Q _07808_/A _07800_/X _07811_/A _07872_/X vssd1 vssd1 vccd1 vccd1
+ _14132_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06826_ _14607_/Q _06823_/X _06825_/X _06811_/X _06821_/X vssd1 vssd1 vccd1 vccd1
+ _14607_/D sky130_fd_sc_hd__o221a_1
X_09614_ _06897_/X _09613_/X _06897_/X _09613_/X vssd1 vssd1 vccd1 vccd1 _09614_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _09545_/A vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06757_ _08126_/A vssd1 vssd1 vccd1 vccd1 _06757_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09476_ _13279_/Q _09472_/X _12274_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _13279_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ _06603_/Y _08962_/A _08957_/A _06628_/Y vssd1 vssd1 vccd1 vccd1 _06688_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08427_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08427_/X sky130_fd_sc_hd__clkbuf_2
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _13890_/Q _08354_/X _08114_/X _08356_/X _08349_/X vssd1 vssd1 vccd1 vccd1
+ _13890_/D sky130_fd_sc_hd__o221a_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07309_ _07309_/A vssd1 vssd1 vccd1 vccd1 _07309_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08289_ _13929_/Q _08284_/X _08114_/X _08286_/X _08288_/X vssd1 vssd1 vccd1 vccd1
+ _13929_/D sky130_fd_sc_hd__o221a_1
XFILLER_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _13193_/Q _10276_/X _14016_/Q _10203_/X _10319_/X vssd1 vssd1 vccd1 vccd1
+ _10320_/X sky130_fd_sc_hd__a221o_2
XFILLER_101_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10251_ _10251_/A vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10182_ _13858_/Q vssd1 vssd1 vccd1 vccd1 _10182_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput590 _13277_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13941_ _14100_/CLK _13941_/D vssd1 vssd1 vccd1 vccd1 _13941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13872_ _14107_/CLK _13872_/D vssd1 vssd1 vccd1 vccd1 _13872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ _12517_/X _12822_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12823_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12754_ _09552_/X _12753_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__mux2_1
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11705_ _11700_/Y _11633_/X _11701_/Y _11635_/X _11704_/X vssd1 vssd1 vccd1 vccd1
+ _11740_/A sky130_fd_sc_hd__o221a_2
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12685_ _09591_/X _12684_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__mux2_1
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _13686_/Q vssd1 vssd1 vccd1 vccd1 _11636_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14424_ _14595_/CLK _14424_/D vssd1 vssd1 vccd1 vccd1 _14424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _14629_/CLK _14355_/D vssd1 vssd1 vccd1 vccd1 _14355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11567_ _11565_/Y _11424_/X _11566_/Y _11426_/X vssd1 vssd1 vccd1 vccd1 _11567_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10518_ _10475_/X _10518_/B _10518_/C _10518_/D vssd1 vssd1 vccd1 vccd1 _10519_/D
+ sky130_fd_sc_hd__and4b_1
X_13306_ _13370_/CLK _13306_/D vssd1 vssd1 vccd1 vccd1 _13306_/Q sky130_fd_sc_hd__dfxtp_1
X_14286_ _14325_/CLK _14286_/D vssd1 vssd1 vccd1 vccd1 _14286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11498_ _11496_/Y _11449_/X _11497_/Y _11451_/X vssd1 vssd1 vccd1 vccd1 _11498_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13237_ _13368_/CLK _13237_/D vssd1 vssd1 vccd1 vccd1 _13269_/Q sky130_fd_sc_hd__dfxtp_2
X_10449_ _13863_/Q vssd1 vssd1 vccd1 vccd1 _10449_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _12663_/X input348/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13168_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12119_ vssd1 vssd1 vccd1 vccd1 _12119_/HI _12119_/LO sky130_fd_sc_hd__conb_1
XFILLER_135_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13099_ _12627_/X _13098_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07660_ _14233_/Q _07653_/X _07345_/X _07654_/X _07658_/X vssd1 vssd1 vccd1 vccd1
+ _14233_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06611_ _06611_/A vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07591_ _14271_/Q _07589_/X _07349_/X _07590_/X _07585_/X vssd1 vssd1 vccd1 vccd1
+ _14271_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09330_ _09519_/A vssd1 vssd1 vccd1 vccd1 _09330_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06542_ _06538_/Y _08825_/A _08822_/A _06541_/Y vssd1 vssd1 vccd1 vccd1 _06542_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09261_ _13429_/Q _09257_/X _09051_/X _09258_/X _09260_/X vssd1 vssd1 vccd1 vccd1
+ _13429_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08212_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08247_/A sky130_fd_sc_hd__buf_4
XFILLER_163_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09192_ _13468_/Q _09188_/X _09051_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1
+ _13468_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08143_ _13996_/Q _08136_/X _08142_/X _08138_/X _08134_/X vssd1 vssd1 vccd1 vccd1
+ _13996_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08074_ _08133_/A vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_159_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07025_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput307 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _06493_/C sky130_fd_sc_hd__clkbuf_1
XPHY_7328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput318 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 _06496_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08976_ _13584_/Q _08969_/X _08974_/X _08971_/X _08975_/X vssd1 vssd1 vccd1 vccd1
+ _13584_/D sky130_fd_sc_hd__o221a_1
Xinput329 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _06488_/B sky130_fd_sc_hd__clkbuf_2
XPHY_6605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07927_ _07927_/A vssd1 vssd1 vccd1 vccd1 _07927_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07858_ _14144_/Q _07855_/X _07771_/X _07856_/X _07857_/X vssd1 vssd1 vccd1 vccd1
+ _14144_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06809_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07789_ _14176_/Q _07783_/X _07788_/X _07785_/X _07781_/X vssd1 vssd1 vccd1 vccd1
+ _14176_/D sky130_fd_sc_hd__o221a_1
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09528_ _09533_/A _12412_/X vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__and2_1
XFILLER_73_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09459_ _09603_/A _09604_/A vssd1 vssd1 vccd1 vccd1 _09459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _12509_/X _06946_/Y _12470_/S vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14140_ _14143_/CLK _14140_/D vssd1 vssd1 vccd1 vccd1 _14140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11352_ _11347_/Y _11219_/X _11348_/Y _11221_/X _11351_/X vssd1 vssd1 vccd1 vccd1
+ _11353_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _10301_/Y _10156_/X _10302_/Y _10159_/X vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14071_ _14071_/CLK _14071_/D vssd1 vssd1 vccd1 vccd1 _14071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11283_ _13880_/Q vssd1 vssd1 vccd1 vccd1 _11283_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13022_ _13021_/X _12590_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13022_/X sky130_fd_sc_hd__mux2_1
X_10234_ _10234_/A vssd1 vssd1 vccd1 vccd1 _10234_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10165_ _10165_/A vssd1 vssd1 vccd1 vccd1 _11831_/A sky130_fd_sc_hd__inv_2
XFILLER_117_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10096_ _10099_/A _10136_/A vssd1 vssd1 vccd1 vccd1 _12476_/S sky130_fd_sc_hd__or2_1
XFILLER_208_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13924_ _14119_/CLK _13924_/D vssd1 vssd1 vccd1 vccd1 _13924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13855_ _14095_/CLK _13855_/D vssd1 vssd1 vccd1 vccd1 _13855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12806_ _12513_/X _12805_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13786_ _14121_/CLK _13786_/D vssd1 vssd1 vccd1 vccd1 _13786_/Q sky130_fd_sc_hd__dfxtp_1
X_10998_ _10996_/Y _10927_/X _10997_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _10998_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12737_ _09541_/X _12736_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12737_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ _09580_/X input359/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__mux2_1
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _14481_/CLK _14407_/D vssd1 vssd1 vccd1 vccd1 _14407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11619_ _13607_/Q vssd1 vssd1 vccd1 vccd1 _11619_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12599_ _09914_/Y _13313_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12599_/X sky130_fd_sc_hd__mux2_1
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14611_/CLK _14338_/D vssd1 vssd1 vccd1 vccd1 _14338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14269_ _14495_/CLK _14269_/D vssd1 vssd1 vccd1 vccd1 _14269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08830_ _13651_/Q _08818_/X _08829_/X _08820_/X _08823_/X vssd1 vssd1 vccd1 vccd1
+ _13651_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08761_ _08777_/A vssd1 vssd1 vccd1 vccd1 _08761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07712_ _07712_/A vssd1 vssd1 vccd1 vccd1 _07712_/X sky130_fd_sc_hd__buf_4
XFILLER_26_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08692_ _13726_/Q _08687_/X _08606_/X _08689_/X _08684_/X vssd1 vssd1 vccd1 vccd1
+ _13726_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07643_ _07687_/A vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__buf_4
XFILLER_4_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07574_ _14281_/Q _07571_/X _07323_/X _07573_/X _07566_/X vssd1 vssd1 vccd1 vccd1
+ _14281_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _13400_/Q _09310_/X _08153_/A _09311_/X _09306_/X vssd1 vssd1 vccd1 vccd1
+ _13400_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06525_ _08989_/D vssd1 vssd1 vccd1 vccd1 _09271_/D sky130_fd_sc_hd__buf_1
XFILLER_39_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09244_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09244_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09175_ _13478_/Q _09171_/X _08948_/X _09172_/X _09173_/X vssd1 vssd1 vccd1 vccd1
+ _13478_/D sky130_fd_sc_hd__o221a_1
XFILLER_182_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08126_ _08126_/A vssd1 vssd1 vccd1 vccd1 _08126_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_198_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08057_ _14035_/Q _08053_/X _07751_/X _08054_/X _08050_/X vssd1 vssd1 vccd1 vccd1
+ _14035_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07008_ _09131_/C vssd1 vssd1 vccd1 vccd1 _08814_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_89_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput104 la_data_in[43] vssd1 vssd1 vccd1 vccd1 _06657_/A sky130_fd_sc_hd__buf_2
XPHY_7125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput115 la_data_in[53] vssd1 vssd1 vccd1 vccd1 _06696_/A sky130_fd_sc_hd__clkbuf_4
XPHY_7136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput126 la_data_in[63] vssd1 vssd1 vccd1 vccd1 _06540_/A sky130_fd_sc_hd__buf_2
XPHY_7147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput137 la_data_in[73] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__buf_1
XPHY_7158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput148 la_data_in[83] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_1
XPHY_7169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput159 la_data_in[93] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__buf_1
X_08959_ _13591_/Q _08956_/X _08957_/X _08958_/X _08951_/X vssd1 vssd1 vccd1 vccd1
+ _13591_/D sky130_fd_sc_hd__o221a_1
XPHY_6435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _14519_/Q vssd1 vssd1 vccd1 vccd1 _11970_/Y sky130_fd_sc_hd__inv_2
XPHY_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10921_ _10921_/A _10921_/B _10921_/C _10921_/D vssd1 vssd1 vccd1 vccd1 _10921_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _13832_/Q vssd1 vssd1 vccd1 vccd1 _10852_/Y sky130_fd_sc_hd__inv_2
X_13640_ _14146_/CLK _13640_/D vssd1 vssd1 vccd1 vccd1 _13640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _14123_/CLK _13571_/D vssd1 vssd1 vccd1 vccd1 _13571_/Q sky130_fd_sc_hd__dfxtp_1
X_10783_ _10778_/Y _10725_/X _10779_/Y _10727_/X _10782_/X vssd1 vssd1 vccd1 vccd1
+ _10796_/B sky130_fd_sc_hd__o221a_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12522_ _13362_/Q _10041_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12522_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12453_ _12452_/X _06924_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12453_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11404_ _11400_/Y _11401_/X _11402_/Y _11403_/X vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__o22a_2
X_12384_ _13210_/Q _12383_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14123_ _14123_/CLK _14123_/D vssd1 vssd1 vccd1 vccd1 _14123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11335_ _14505_/Q vssd1 vssd1 vccd1 vccd1 _11335_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14054_ _14056_/CLK _14054_/D vssd1 vssd1 vccd1 vccd1 _14054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11266_ _13482_/Q vssd1 vssd1 vccd1 vccd1 _11266_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10217_ _10217_/A vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__clkbuf_2
X_13005_ _12582_/X _13004_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11197_ _13211_/Q _11013_/X _14034_/Q _11193_/X _11196_/X vssd1 vssd1 vccd1 vccd1
+ _11197_/X sky130_fd_sc_hd__a221o_4
XFILLER_171_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10148_ _14053_/Q vssd1 vssd1 vccd1 vccd1 _10148_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ _10079_/A _10125_/A vssd1 vssd1 vccd1 vccd1 _12491_/S sky130_fd_sc_hd__or2_1
XFILLER_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13907_ _14143_/CLK _13907_/D vssd1 vssd1 vccd1 vccd1 _13907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13838_ _13996_/CLK _13838_/D vssd1 vssd1 vccd1 vccd1 _13838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _14120_/CLK _13769_/D vssd1 vssd1 vccd1 vccd1 _13769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07290_ _07290_/A vssd1 vssd1 vccd1 vccd1 _07290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09931_ _09931_/A vssd1 vssd1 vccd1 vccd1 _09931_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09862_ _13306_/Q vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__inv_2
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08813_ _08813_/A vssd1 vssd1 vccd1 vccd1 _09132_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_154_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__or2_1
XFILLER_45_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _08744_/A _09201_/B _08744_/C _09201_/D vssd1 vssd1 vccd1 vccd1 _11637_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08675_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__inv_2
XPHY_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_209 _13279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07626_ _14248_/Q _07561_/A _07480_/X _07563_/A _07624_/X vssd1 vssd1 vccd1 vccd1
+ _14248_/D sky130_fd_sc_hd__o221a_1
XPHY_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ _09271_/A _09063_/B _09131_/C _08673_/D vssd1 vssd1 vccd1 vccd1 _11685_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06508_ _06508_/A _06508_/B vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__or2_1
XFILLER_39_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07488_ _07488_/A vssd1 vssd1 vccd1 vccd1 _07488_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09227_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__buf_2
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _13489_/Q _09155_/X _08917_/X _09156_/X _09157_/X vssd1 vssd1 vccd1 vccd1
+ _13489_/D sky130_fd_sc_hd__o221a_1
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08109_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08109_/X sky130_fd_sc_hd__clkbuf_2
X_09089_ _13527_/Q _09086_/X _08920_/X _09087_/X _09084_/X vssd1 vssd1 vccd1 vccd1
+ _13527_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _13441_/Q vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ _11049_/Y _10947_/X _11050_/Y _10949_/X vssd1 vssd1 vccd1 vccd1 _11051_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_192_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10002_ _13372_/Q _10002_/B vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__nand2_4
XFILLER_24_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _11951_/Y _10156_/A _11952_/Y _10159_/A vssd1 vssd1 vccd1 vccd1 _11953_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_6298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ _14613_/Q vssd1 vssd1 vccd1 vccd1 _10904_/Y sky130_fd_sc_hd__inv_2
XPHY_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _11882_/Y _10195_/A _11883_/Y _10198_/A vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ _14047_/CLK _13623_/D vssd1 vssd1 vccd1 vccd1 _13623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10835_ _14455_/Q vssd1 vssd1 vccd1 vccd1 _10835_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _14114_/CLK _13554_/D vssd1 vssd1 vccd1 vccd1 _13554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10766_ _13869_/Q vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12505_ _12504_/X _06996_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12505_/X sky130_fd_sc_hd__mux2_2
XFILLER_199_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10697_ _10697_/A vssd1 vssd1 vccd1 vccd1 _10697_/X sky130_fd_sc_hd__clkbuf_4
X_13485_ _14470_/CLK _13485_/D vssd1 vssd1 vccd1 vccd1 _13485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ _12435_/X _06902_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput408 _12087_/LO vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput419 _12235_/A vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12367_ _12366_/X _13200_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12367_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ _14110_/CLK _14106_/D vssd1 vssd1 vccd1 vccd1 _14106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11318_ _11316_/Y _11165_/X _11317_/Y _11167_/X vssd1 vssd1 vccd1 vccd1 _11318_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_64_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12298_ _11395_/Y _14545_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12298_/X sky130_fd_sc_hd__mux2_2
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11249_ _11485_/A vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__buf_4
X_14037_ _14114_/CLK _14037_/D vssd1 vssd1 vccd1 vccd1 _14037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06790_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08460_ _08460_/A vssd1 vssd1 vccd1 vccd1 _08460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07411_ _07411_/A vssd1 vssd1 vccd1 vccd1 _07411_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08391_ _13870_/Q _08388_/X _08165_/X _08389_/X _08384_/X vssd1 vssd1 vccd1 vccd1
+ _13870_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07342_ _14391_/Q _07335_/X _07341_/X _07337_/X _07333_/X vssd1 vssd1 vccd1 vccd1
+ _14391_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07273_ _14423_/Q _07265_/X _06784_/X _07266_/X _07271_/X vssd1 vssd1 vccd1 vccd1
+ _14423_/D sky130_fd_sc_hd__o221a_1
X_09012_ _13569_/Q _09004_/X _08912_/X _09006_/X _09011_/X vssd1 vssd1 vccd1 vccd1
+ _13569_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _09912_/A _09912_/B _09913_/Y vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09845_ _13334_/Q _09843_/Y _09785_/B vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09776_ _09776_/A _09776_/B vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__or2_1
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06988_ _14564_/Q vssd1 vssd1 vccd1 vccd1 _06989_/A sky130_fd_sc_hd__inv_2
XFILLER_2_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _13705_/Q _08722_/X _08560_/X _08723_/X _08720_/X vssd1 vssd1 vccd1 vccd1
+ _13705_/D sky130_fd_sc_hd__o221a_1
XPHY_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08658_ _13741_/Q _08588_/A _08657_/X _08591_/A _08653_/X vssd1 vssd1 vccd1 vccd1
+ _13741_/D sky130_fd_sc_hd__o221a_1
XFILLER_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07609_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08895_/A vssd1 vssd1 vccd1 vccd1 _08589_/X sky130_fd_sc_hd__buf_2
XFILLER_109_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10620_ _13508_/Q vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__inv_2
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10551_ _14254_/Q vssd1 vssd1 vccd1 vccd1 _10551_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10482_ _14604_/Q vssd1 vssd1 vccd1 vccd1 _10482_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13270_ _13877_/CLK _13270_/D vssd1 vssd1 vccd1 vccd1 _13270_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ vssd1 vssd1 vccd1 vccd1 _12152_/HI _12152_/LO sky130_fd_sc_hd__conb_1
XFILLER_159_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11103_ _11101_/Y _10967_/X _11102_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _11103_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12083_ vssd1 vssd1 vccd1 vccd1 _12083_/HI _12083_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11034_ _11015_/X _11034_/B _11034_/C _11034_/D vssd1 vssd1 vccd1 vccd1 _11035_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _12572_/X _12984_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _12985_/X sky130_fd_sc_hd__mux2_1
XPHY_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11936_ _13614_/Q vssd1 vssd1 vccd1 vccd1 _11936_/Y sky130_fd_sc_hd__inv_2
XPHY_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _14088_/Q vssd1 vssd1 vccd1 vccd1 _11867_/Y sky130_fd_sc_hd__inv_2
XPHY_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13606_ _14529_/CLK _13606_/D vssd1 vssd1 vccd1 vccd1 _13606_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10818_ _13551_/Q _10720_/X _13792_/Q _10721_/X vssd1 vssd1 vccd1 vccd1 _10818_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14586_ _14621_/CLK _14586_/D vssd1 vssd1 vccd1 vccd1 _14586_/Q sky130_fd_sc_hd__dfxtp_1
X_11798_ _14008_/Q vssd1 vssd1 vccd1 vccd1 _11798_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13537_ _14130_/CLK _13537_/D vssd1 vssd1 vccd1 vccd1 _13537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _11459_/A vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13468_ _14178_/CLK _13468_/D vssd1 vssd1 vccd1 vccd1 _13468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12419_ _12509_/X _06875_/Y _12419_/S vssd1 vssd1 vccd1 vccd1 _12419_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13399_ _14188_/CLK _13399_/D vssd1 vssd1 vccd1 vccd1 _13399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07960_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06911_ _06917_/A _06911_/B vssd1 vssd1 vccd1 vccd1 _14586_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07891_ _07934_/A vssd1 vssd1 vccd1 vccd1 _07926_/A sky130_fd_sc_hd__buf_4
XFILLER_68_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09630_ _14595_/Q _14590_/Q _06872_/Y _06893_/X vssd1 vssd1 vccd1 vccd1 _09630_/X
+ sky130_fd_sc_hd__o22a_1
X_06842_ _08981_/A vssd1 vssd1 vccd1 vccd1 _06843_/B sky130_fd_sc_hd__buf_8
XFILLER_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09561_ _09557_/X _09560_/X _13270_/Q _09558_/X vssd1 vssd1 vccd1 vccd1 _13238_/D
+ sky130_fd_sc_hd__o22a_1
X_06773_ _14622_/Q _06769_/X _06771_/X _06772_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _14622_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08512_ _13809_/Q _08500_/X _08510_/X _08503_/X _08511_/X vssd1 vssd1 vccd1 vccd1
+ _13809_/D sky130_fd_sc_hd__o221a_1
XFILLER_188_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09492_ _13267_/Q _09486_/X _12262_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _13267_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ _13843_/Q _08436_/X _08132_/X _08437_/X _08441_/X vssd1 vssd1 vccd1 vccd1
+ _13843_/D sky130_fd_sc_hd__o221a_1
XFILLER_93_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _13880_/Q _08371_/X _08140_/X _08372_/X _08367_/X vssd1 vssd1 vccd1 vccd1
+ _13880_/D sky130_fd_sc_hd__o221a_1
XFILLER_205_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07325_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07325_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07256_ _14433_/Q _07248_/X _06748_/X _07250_/X _07254_/X vssd1 vssd1 vccd1 vccd1
+ _14433_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _14471_/Q _07185_/X _06753_/X _07186_/X _07181_/X vssd1 vssd1 vccd1 vccd1
+ _14471_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09828_ _09789_/A _09789_/B _09827_/Y vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09759_ _13329_/Q vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__inv_2
XFILLER_55_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12770_ _09519_/X _12769_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__mux2_1
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _14513_/Q vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__inv_2
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14440_ _14481_/CLK _14440_/D vssd1 vssd1 vccd1 vccd1 _14440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11652_ _13849_/Q vssd1 vssd1 vccd1 vccd1 _11652_/Y sky130_fd_sc_hd__inv_2
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10603_ _10603_/A _10603_/B _10603_/C _10603_/D vssd1 vssd1 vccd1 vccd1 _10603_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14371_ _14629_/CLK _14371_/D vssd1 vssd1 vccd1 vccd1 _14371_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11583_ _13925_/Q vssd1 vssd1 vccd1 vccd1 _11583_/Y sky130_fd_sc_hd__inv_2
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _13352_/CLK _13322_/D vssd1 vssd1 vccd1 vccd1 _13322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534_ _10532_/Y _10455_/X _10533_/Y _10458_/X vssd1 vssd1 vccd1 vccd1 _10534_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10465_ _11426_/A vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13253_ _13372_/CLK _13253_/D vssd1 vssd1 vccd1 vccd1 _13285_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12204_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10396_ _10394_/Y _10188_/X _10395_/Y _10191_/X vssd1 vssd1 vccd1 vccd1 _10396_/X
+ sky130_fd_sc_hd__o22a_1
X_13184_ _13180_/X _13181_/X _13182_/X _13183_/X _12510_/S _10058_/B vssd1 vssd1 vccd1
+ vccd1 _13184_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ vssd1 vssd1 vccd1 vccd1 _12135_/HI _12135_/LO sky130_fd_sc_hd__conb_1
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12066_ _09793_/A _12064_/X _09905_/A _12065_/X vssd1 vssd1 vccd1 vccd1 _12066_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11017_ _14342_/Q vssd1 vssd1 vccd1 vccd1 _11017_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _12564_/X input333/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__mux2_1
XPHY_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11919_ _11917_/Y _10181_/A _11918_/Y _10184_/A vssd1 vssd1 vccd1 vccd1 _11919_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12535_/X _12898_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12899_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14638_ _14639_/CLK _14638_/D vssd1 vssd1 vccd1 vccd1 _14639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14569_ _14573_/CLK _14569_/D vssd1 vssd1 vccd1 vccd1 _14569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07110_ _14511_/Q _07102_/X _06748_/X _07104_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _14511_/D sky130_fd_sc_hd__o221a_1
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ _14014_/Q _08025_/A _07876_/X _08027_/A _08089_/X vssd1 vssd1 vccd1 vccd1
+ _14014_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07041_ _14547_/Q _07035_/X _06760_/X _07036_/X _07038_/X vssd1 vssd1 vccd1 vccd1
+ _14547_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _09048_/A vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07943_ _14097_/Q _07934_/X _07790_/X _07935_/X _07940_/X vssd1 vssd1 vccd1 vccd1
+ _14097_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07874_ _14133_/Q _07808_/A _07798_/X _07811_/A _07872_/X vssd1 vssd1 vccd1 vccd1
+ _14133_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09613_ _06961_/Y _14568_/Q _14572_/Q _06975_/Y vssd1 vssd1 vccd1 vccd1 _09613_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06825_ _08175_/A vssd1 vssd1 vccd1 vccd1 _06825_/X sky130_fd_sc_hd__buf_2
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09544_ _09557_/A vssd1 vssd1 vccd1 vccd1 _09544_/X sky130_fd_sc_hd__clkbuf_2
X_06756_ _08920_/A vssd1 vssd1 vccd1 vccd1 _08126_/A sky130_fd_sc_hd__buf_4
XFILLER_37_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ _13280_/Q _09472_/X _12275_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _13280_/D
+ sky130_fd_sc_hd__o22a_1
X_06687_ _06678_/X _06686_/X _06678_/X _06686_/X vssd1 vssd1 vccd1 vccd1 _06853_/B
+ sky130_fd_sc_hd__a2bb2o_2
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08426_ _08469_/A vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08357_ _13891_/Q _08354_/X _08110_/X _08356_/X _08349_/X vssd1 vssd1 vccd1 vccd1
+ _13891_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07308_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08288_ _08288_/A vssd1 vssd1 vccd1 vccd1 _08288_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07239_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10250_ _11695_/A vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput580 _13268_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput591 _13278_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _14100_/CLK _13940_/D vssd1 vssd1 vccd1 vccd1 _13940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _14107_/CLK _13871_/D vssd1 vssd1 vccd1 vccd1 _13871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12822_ _12517_/X _12821_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12822_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ _09552_/X _12752_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12753_/X sky130_fd_sc_hd__mux2_1
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11704_ _11702_/Y _11637_/X _11703_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _11704_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12684_ _09591_/X input355/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__mux2_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14423_ _14573_/CLK _14423_/D vssd1 vssd1 vccd1 vccd1 _14423_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11635_ _11635_/A vssd1 vssd1 vccd1 vccd1 _11635_/X sky130_fd_sc_hd__buf_2
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14354_ _14629_/CLK _14354_/D vssd1 vssd1 vccd1 vccd1 _14354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _13528_/Q vssd1 vssd1 vccd1 vccd1 _11566_/Y sky130_fd_sc_hd__inv_2
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13305_ _13368_/CLK _13305_/D vssd1 vssd1 vccd1 vccd1 _13305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10517_ _10504_/Y _10506_/X _10507_/Y _10509_/X _10516_/X vssd1 vssd1 vccd1 vccd1
+ _10518_/D sky130_fd_sc_hd__o221a_1
X_14285_ _14325_/CLK _14285_/D vssd1 vssd1 vccd1 vccd1 _14285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11497_ _14274_/Q vssd1 vssd1 vccd1 vccd1 _11497_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _13352_/CLK _13236_/D vssd1 vssd1 vccd1 vccd1 _13268_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _11414_/A vssd1 vssd1 vccd1 vccd1 _10448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13167_ _12661_/X _13166_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10379_ _10374_/Y _10242_/X _10375_/Y _10245_/X _10378_/X vssd1 vssd1 vccd1 vccd1
+ _10380_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12118_ vssd1 vssd1 vccd1 vccd1 _12118_/HI _12118_/LO sky130_fd_sc_hd__conb_1
X_13098_ _13097_/X _12627_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12049_ _09782_/A _12043_/X _09894_/A _12044_/X vssd1 vssd1 vccd1 vccd1 _12049_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06610_ _06582_/Y _08940_/A _08933_/A _06554_/Y vssd1 vssd1 vccd1 vccd1 _06699_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07590_ _07606_/A vssd1 vssd1 vccd1 vccd1 _07590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06541_ _06541_/A vssd1 vssd1 vccd1 vccd1 _06541_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09260_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08211_ _08246_/A vssd1 vssd1 vccd1 vccd1 _08211_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ _13469_/Q _09188_/X _08970_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1
+ _13469_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08142_ _08142_/A vssd1 vssd1 vccd1 vccd1 _08142_/X sky130_fd_sc_hd__buf_4
XFILLER_198_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08073_ _14025_/Q _08069_/X _07776_/X _08070_/X _08066_/X vssd1 vssd1 vccd1 vccd1
+ _14025_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__buf_4
XFILLER_192_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput308 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _06499_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08975_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08975_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput319 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _06512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07926_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07926_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07857_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06808_ _14612_/Q _06805_/X _06807_/X _06790_/X _06803_/X vssd1 vssd1 vccd1 vccd1
+ _14612_/D sky130_fd_sc_hd__o221a_1
X_07788_ _08179_/A vssd1 vssd1 vccd1 vccd1 _07788_/X sky130_fd_sc_hd__buf_4
XFILLER_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _09514_/X _09526_/X _13282_/Q _09517_/X vssd1 vssd1 vccd1 vccd1 _13250_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06739_ _14631_/Q _06733_/X _06738_/X _06726_/X _06730_/X vssd1 vssd1 vccd1 vccd1
+ _14631_/D sky130_fd_sc_hd__o221a_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09458_/A _12262_/S vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__or2_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08409_ _08813_/A vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__buf_2
XFILLER_36_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09389_ _09509_/A vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__buf_4
XFILLER_200_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _14117_/Q vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _11349_/Y _11223_/X _11350_/Y _11225_/X vssd1 vssd1 vccd1 vccd1 _11351_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _13619_/Q vssd1 vssd1 vccd1 vccd1 _10302_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14070_ _14071_/CLK _14070_/D vssd1 vssd1 vccd1 vccd1 _14070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11282_ _13763_/Q vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _12590_/X _13020_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__mux2_1
X_10233_ _11683_/A vssd1 vssd1 vccd1 vccd1 _10234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _10696_/A vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10095_ _10107_/B _10132_/A vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__or2_1
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13923_ _14119_/CLK _13923_/D vssd1 vssd1 vccd1 vccd1 _13923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _14095_/CLK _13854_/D vssd1 vssd1 vccd1 vccd1 _13854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12805_ _12513_/X _12804_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13785_ _14121_/CLK _13785_/D vssd1 vssd1 vccd1 vccd1 _13785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10997_ _13633_/Q vssd1 vssd1 vccd1 vccd1 _10997_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12736_ _09541_/X input344/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12736_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _13343_/Q _12666_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__mux2_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _14481_/CLK _14406_/D vssd1 vssd1 vccd1 vccd1 _14406_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11618_ _14316_/Q vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12598_ _13314_/Q _12597_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__mux2_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14337_ _14611_/CLK _14337_/D vssd1 vssd1 vccd1 vccd1 _14337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11549_ _11549_/A _11549_/B _11549_/C _11549_/D vssd1 vssd1 vccd1 vccd1 _11549_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_7_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14268_ _14495_/CLK _14268_/D vssd1 vssd1 vccd1 vccd1 _14268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13219_ _13350_/CLK _13219_/D vssd1 vssd1 vccd1 vccd1 _13219_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14199_ _14291_/CLK _14199_/D vssd1 vssd1 vccd1 vccd1 _14199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08760_ _08793_/A vssd1 vssd1 vccd1 vccd1 _08760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07711_ _14206_/Q _07704_/X _07710_/X _07706_/X _07698_/X vssd1 vssd1 vccd1 vccd1
+ _14206_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08691_ _13727_/Q _08687_/X _08505_/X _08689_/X _08684_/X vssd1 vssd1 vccd1 vccd1
+ _13727_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07642_ _14243_/Q _07634_/X _07317_/X _07636_/X _07640_/X vssd1 vssd1 vccd1 vccd1
+ _14243_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07573_ _07606_/A vssd1 vssd1 vccd1 vccd1 _07573_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09312_ _13401_/Q _09310_/X _08150_/A _09311_/X _09306_/X vssd1 vssd1 vccd1 vccd1
+ _13401_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06524_ input89/X _07232_/B vssd1 vssd1 vccd1 vccd1 _08989_/C sky130_fd_sc_hd__or2_2
XFILLER_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09243_ _13440_/Q _09241_/X _08945_/X _09242_/X _09236_/X vssd1 vssd1 vccd1 vccd1
+ _13440_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09174_ _13479_/Q _09171_/X _08945_/X _09172_/X _09173_/X vssd1 vssd1 vccd1 vccd1
+ _13479_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08125_ _14003_/Q _08122_/X _08123_/X _08124_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _14003_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ _14036_/Q _08053_/X _07749_/X _08054_/X _08050_/X vssd1 vssd1 vccd1 vccd1
+ _14036_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07007_ input89/X _07086_/B vssd1 vssd1 vccd1 vccd1 _09131_/C sky130_fd_sc_hd__or2_2
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput105 la_data_in[44] vssd1 vssd1 vccd1 vccd1 _06602_/A sky130_fd_sc_hd__buf_2
XPHY_7126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 la_data_in[54] vssd1 vssd1 vccd1 vccd1 _06626_/A sky130_fd_sc_hd__buf_2
XPHY_7137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 la_data_in[64] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
XPHY_7148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput138 la_data_in[74] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__buf_1
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08958_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__clkbuf_2
XPHY_7159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput149 la_data_in[84] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__buf_1
XFILLER_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ _14116_/Q _07902_/X _07742_/X _07903_/X _07905_/X vssd1 vssd1 vccd1 vccd1
+ _14116_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _13617_/Q _08818_/A _08657_/X _08820_/A _08886_/X vssd1 vssd1 vccd1 vccd1
+ _13617_/D sky130_fd_sc_hd__o221a_1
XPHY_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _10901_/X _10920_/B _10920_/C _10920_/D vssd1 vssd1 vccd1 vccd1 _10921_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _10849_/Y _10704_/X _10850_/Y _10706_/X vssd1 vssd1 vccd1 vccd1 _10851_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _14121_/CLK _13570_/D vssd1 vssd1 vccd1 vccd1 _13570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10782_ _10780_/Y _10729_/X _10781_/Y _10731_/X vssd1 vssd1 vccd1 vccd1 _10782_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12521_ _13363_/Q _10042_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__mux2_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12452_ _12509_/X _06924_/Y _12452_/S vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _11403_/A vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12383_ _13210_/Q _06614_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14122_ _14123_/CLK _14122_/D vssd1 vssd1 vccd1 vccd1 _14122_/Q sky130_fd_sc_hd__dfxtp_1
X_11334_ _13214_/Q _11249_/X _14037_/Q _11193_/X _11333_/X vssd1 vssd1 vccd1 vccd1
+ _11334_/X sky130_fd_sc_hd__a221o_4
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14053_ _14056_/CLK _14053_/D vssd1 vssd1 vccd1 vccd1 _14053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11265_ _14152_/Q vssd1 vssd1 vccd1 vccd1 _11265_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _12582_/X input340/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10216_ _11671_/A vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__buf_2
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11196_ _13559_/Q _11194_/X _13800_/Q _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10147_ _10147_/A vssd1 vssd1 vccd1 vccd1 _12322_/S sky130_fd_sc_hd__clkinv_8
XFILLER_153_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10078_ _10102_/B _10122_/A vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__or2_1
XFILLER_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ _14143_/CLK _13906_/D vssd1 vssd1 vccd1 vccd1 _13906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13837_ _14107_/CLK _13837_/D vssd1 vssd1 vccd1 vccd1 _13837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13768_ _14120_/CLK _13768_/D vssd1 vssd1 vccd1 vccd1 _13768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12719_ _09569_/X _12718_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13202_/D sky130_fd_sc_hd__mux2_1
X_13699_ _14178_/CLK _13699_/D vssd1 vssd1 vccd1 vccd1 _13699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09930_ _13318_/Q _09927_/Y _09929_/Y _09927_/A vssd1 vssd1 vccd1 vccd1 _09930_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09861_ _13307_/Q vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__inv_2
XFILLER_140_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08812_ _13656_/Q _08748_/A _08657_/X _08750_/A _08808_/X vssd1 vssd1 vccd1 vccd1
+ _13656_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09792_ _09792_/A _09830_/A vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__or2_2
XFILLER_80_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08989_/D vssd1 vssd1 vccd1 vccd1 _09201_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08674_ _08745_/A _10171_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__or2_4
XPHY_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _14249_/Q _07561_/A _07403_/X _07563_/A _07624_/X vssd1 vssd1 vccd1 vccd1
+ _14249_/D sky130_fd_sc_hd__o221a_1
XPHY_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07556_ _08482_/D vssd1 vssd1 vccd1 vccd1 _08673_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06507_ _06507_/A _06507_/B _06507_/C _06507_/D vssd1 vssd1 vccd1 vccd1 _06508_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_35_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07487_ _07541_/A vssd1 vssd1 vccd1 vccd1 _07488_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _13450_/Q _09224_/X _08917_/X _09225_/X _09219_/X vssd1 vssd1 vccd1 vccd1
+ _13450_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09157_ _09173_/A vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _08174_/A vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__buf_4
XFILLER_11_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09088_ _13528_/Q _09086_/X _08917_/X _09087_/X _09084_/X vssd1 vssd1 vccd1 vccd1
+ _13528_/D sky130_fd_sc_hd__o221a_1
X_08039_ _14047_/Q _08036_/X _07719_/X _08038_/X _08032_/X vssd1 vssd1 vccd1 vccd1
+ _14047_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11050_ _14109_/Q vssd1 vssd1 vccd1 vccd1 _11050_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10001_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10002_/B sky130_fd_sc_hd__inv_2
XFILLER_133_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _13654_/Q vssd1 vssd1 vccd1 vccd1 _11952_/Y sky130_fd_sc_hd__inv_2
XPHY_6288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10903_ _14340_/Q vssd1 vssd1 vccd1 vccd1 _10903_/Y sky130_fd_sc_hd__inv_2
XPHY_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11883_ _13535_/Q vssd1 vssd1 vccd1 vccd1 _11883_/Y sky130_fd_sc_hd__inv_2
XPHY_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ _14047_/CLK _13622_/D vssd1 vssd1 vccd1 vccd1 _13622_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ _13473_/Q vssd1 vssd1 vccd1 vccd1 _10834_/Y sky130_fd_sc_hd__inv_2
XPHY_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _14114_/CLK _13553_/D vssd1 vssd1 vccd1 vccd1 _13553_/Q sky130_fd_sc_hd__dfxtp_1
X_10765_ _13752_/Q vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _12503_/X _06996_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13484_ _14595_/CLK _13484_/D vssd1 vssd1 vccd1 vccd1 _13484_/Q sky130_fd_sc_hd__dfxtp_1
X_10696_ _10696_/A vssd1 vssd1 vccd1 vccd1 _10696_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_199_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _12434_/X _06902_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12435_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12366_ _13200_/Q _12365_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__mux2_1
Xoutput409 _12088_/LO vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _14110_/CLK _14105_/D vssd1 vssd1 vccd1 vccd1 _14105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11317_ _13640_/Q vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _11465_/Y _14546_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12297_/X sky130_fd_sc_hd__mux2_2
XFILLER_113_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14036_ _14114_/CLK _14036_/D vssd1 vssd1 vccd1 vccd1 _14036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11248_ _11238_/Y _11176_/X _11241_/X _11244_/X _11247_/X vssd1 vssd1 vccd1 vccd1
+ _11271_/C sky130_fd_sc_hd__o2111a_4
XFILLER_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _13878_/Q vssd1 vssd1 vccd1 vccd1 _11179_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07410_ _07467_/A vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08390_ _13871_/Q _08388_/X _08162_/X _08389_/X _08384_/X vssd1 vssd1 vccd1 vccd1
+ _13871_/D sky130_fd_sc_hd__o221a_1
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07341_ _08128_/A vssd1 vssd1 vccd1 vccd1 _07341_/X sky130_fd_sc_hd__buf_2
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07272_ _14424_/Q _07265_/X _06781_/X _07266_/X _07271_/X vssd1 vssd1 vccd1 vccd1
+ _14424_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _09036_/A vssd1 vssd1 vccd1 vccd1 _09011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09913_ _09916_/B vssd1 vssd1 vccd1 vccd1 _09913_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09844_ _09783_/A _09783_/B _09843_/Y vssd1 vssd1 vccd1 vccd1 _09844_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09775_ _09775_/A _09853_/A vssd1 vssd1 vccd1 vccd1 _09776_/B sky130_fd_sc_hd__or2_1
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06987_ _06991_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _14565_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08726_ _13706_/Q _08722_/X _08558_/X _08723_/X _08720_/X vssd1 vssd1 vccd1 vccd1
+ _13706_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08657_ _09060_/A vssd1 vssd1 vccd1 vccd1 _08657_/X sky130_fd_sc_hd__clkbuf_4
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _14260_/Q _07605_/X _07377_/X _07606_/X _07601_/X vssd1 vssd1 vccd1 vccd1
+ _14260_/D sky130_fd_sc_hd__o221a_1
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08588_ _08588_/A vssd1 vssd1 vccd1 vccd1 _08588_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07539_ _14297_/Q _07532_/X _07381_/X _07533_/X _07536_/X vssd1 vssd1 vccd1 vccd1
+ _14297_/D sky130_fd_sc_hd__o221a_1
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10550_ _14176_/Q vssd1 vssd1 vccd1 vccd1 _10550_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09219_/A vssd1 vssd1 vccd1 vccd1 _09209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10481_ _11437_/A vssd1 vssd1 vccd1 vccd1 _10481_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12151_ vssd1 vssd1 vccd1 vccd1 _12151_/HI _12151_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _14383_/Q vssd1 vssd1 vccd1 vccd1 _11102_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12082_ vssd1 vssd1 vccd1 vccd1 _12082_/HI _12082_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11033_ _11028_/Y _10983_/X _11029_/Y _10985_/X _11032_/X vssd1 vssd1 vccd1 vccd1
+ _11034_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12984_ _12572_/X input360/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12984_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11935_ _14323_/Q vssd1 vssd1 vccd1 vccd1 _11935_/Y sky130_fd_sc_hd__inv_2
XPHY_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11866_ _11866_/A _11866_/B _11866_/C _11866_/D vssd1 vssd1 vccd1 vccd1 _11866_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_127_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _14529_/CLK _13605_/D vssd1 vssd1 vccd1 vccd1 _13605_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ _10807_/Y _10702_/X _10810_/X _10813_/X _10816_/X vssd1 vssd1 vccd1 vccd1
+ _10839_/C sky130_fd_sc_hd__o2111a_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585_ _14621_/CLK _14585_/D vssd1 vssd1 vccd1 vccd1 _14585_/Q sky130_fd_sc_hd__dfxtp_2
X_11797_ _11795_/Y _11653_/X _11796_/Y _11655_/X vssd1 vssd1 vccd1 vccd1 _11797_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13536_ _14130_/CLK _13536_/D vssd1 vssd1 vccd1 vccd1 _13536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10748_ _13471_/Q vssd1 vssd1 vccd1 vccd1 _10748_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13467_ _14178_/CLK _13467_/D vssd1 vssd1 vccd1 vccd1 _13467_/Q sky130_fd_sc_hd__dfxtp_1
X_10679_ _14140_/Q vssd1 vssd1 vccd1 vccd1 _10679_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12418_ _12417_/X _13215_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13398_ _14188_/CLK _13398_/D vssd1 vssd1 vccd1 vccd1 _13398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12349_ _12348_/X _13206_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12349_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14047_/CLK _14019_/D vssd1 vssd1 vccd1 vccd1 _14019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06910_ _06901_/X _12296_/X _06909_/Y _06903_/X vssd1 vssd1 vccd1 vccd1 _06911_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07890_ _14126_/Q _07882_/X _07714_/X _07884_/X _07886_/X vssd1 vssd1 vccd1 vccd1
+ _14126_/D sky130_fd_sc_hd__o221a_1
XFILLER_155_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06841_ _14602_/Q _06530_/A _06532_/X _08186_/A _06838_/X vssd1 vssd1 vccd1 vccd1
+ _14602_/D sky130_fd_sc_hd__o221a_1
XFILLER_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09560_ _09560_/A _12349_/X vssd1 vssd1 vccd1 vccd1 _09560_/X sky130_fd_sc_hd__and2_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06772_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08511_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__clkbuf_2
X_09491_ _13268_/Q _09486_/X _12263_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _13268_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08442_ _13844_/Q _08436_/X _08130_/X _08437_/X _08441_/X vssd1 vssd1 vccd1 vccd1
+ _13844_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _13881_/Q _08371_/X _08137_/X _08372_/X _08367_/X vssd1 vssd1 vccd1 vccd1
+ _13881_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07324_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ _14434_/Q _07248_/X _06745_/X _07250_/X _07254_/X vssd1 vssd1 vccd1 vccd1
+ _14434_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07186_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07186_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _09827_/A vssd1 vssd1 vccd1 vccd1 _09827_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09758_ _13330_/Q vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__inv_2
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08709_ _13717_/Q _08706_/X _08530_/X _08707_/X _08704_/X vssd1 vssd1 vccd1 vccd1
+ _13717_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09689_ _09671_/A _09688_/X _09671_/A _09688_/X vssd1 vssd1 vccd1 vccd1 _09689_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_199_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _13222_/Q _11013_/A _14045_/Q _11663_/X _11719_/X vssd1 vssd1 vccd1 vccd1
+ _11720_/X sky130_fd_sc_hd__a221o_4
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11651_ _11647_/Y _11648_/X _11649_/Y _11650_/X vssd1 vssd1 vccd1 vccd1 _11651_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10602_ _10583_/X _10602_/B _10602_/C _10602_/D vssd1 vssd1 vccd1 vccd1 _10603_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _14629_/CLK _14370_/D vssd1 vssd1 vccd1 vccd1 _14370_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11582_ _11577_/Y _11445_/X _11578_/Y _11447_/X _11581_/X vssd1 vssd1 vccd1 vccd1
+ _11589_/C sky130_fd_sc_hd__o221a_1
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ _13352_/CLK _13321_/D vssd1 vssd1 vccd1 vccd1 _13321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10533_ _14098_/Q vssd1 vssd1 vccd1 vccd1 _10533_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ _13372_/CLK _13252_/D vssd1 vssd1 vccd1 vccd1 _13284_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_183_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10464_ _11660_/A vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12203_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ _14585_/Q _14586_/Q _14583_/Q _14584_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13183_/X sky130_fd_sc_hd__mux4_1
X_10395_ _14096_/Q vssd1 vssd1 vccd1 vccd1 _10395_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12134_ vssd1 vssd1 vccd1 vccd1 _12134_/HI _12134_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12065_ _12065_/A vssd1 vssd1 vccd1 vccd1 _12065_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11016_ _14498_/Q vssd1 vssd1 vccd1 vccd1 _11016_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12967_ _12562_/X _12966_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__mux2_1
XPHY_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11918_ _13894_/Q vssd1 vssd1 vccd1 vccd1 _11918_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12898_ _12535_/X _12897_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14637_ _14637_/CLK _14637_/D vssd1 vssd1 vccd1 vccd1 _14637_/Q sky130_fd_sc_hd__dfxtp_1
X_11849_ _14633_/Q vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14568_ _14573_/CLK _14568_/D vssd1 vssd1 vccd1 vccd1 _14568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13519_ _14114_/CLK _13519_/D vssd1 vssd1 vccd1 vccd1 _13519_/Q sky130_fd_sc_hd__dfxtp_1
X_14499_ _14621_/CLK _14499_/D vssd1 vssd1 vccd1 vccd1 _14499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07040_ _14548_/Q _07035_/X _06757_/X _07036_/X _07038_/X vssd1 vssd1 vccd1 vccd1
+ _14548_/D sky130_fd_sc_hd__o221a_1
XFILLER_155_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08991_ _09049_/A vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__inv_2
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07942_ _14098_/Q _07934_/X _07788_/X _07935_/X _07940_/X vssd1 vssd1 vccd1 vccd1
+ _14098_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07873_ _14134_/Q _07808_/A _07796_/X _07811_/A _07872_/X vssd1 vssd1 vccd1 vccd1
+ _14134_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09612_ _06858_/Y _14575_/Q _14598_/Q _06949_/Y vssd1 vssd1 vccd1 vccd1 _09612_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06824_ input96/X vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09543_ _09547_/A _12379_/X vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__and2_1
X_06755_ _14627_/Q _06751_/X _06753_/X _06754_/X _06749_/X vssd1 vssd1 vccd1 vccd1
+ _14627_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09474_ _13281_/Q _09472_/X _12276_/X _09473_/X vssd1 vssd1 vccd1 vccd1 _13281_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06686_ _06683_/X _06685_/X _06683_/X _06685_/X vssd1 vssd1 vccd1 vccd1 _06686_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08425_ _08460_/A vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__clkbuf_2
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _08389_/A vssd1 vssd1 vccd1 vccd1 _08356_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07307_ _07307_/A vssd1 vssd1 vccd1 vccd1 _07307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08287_ _13930_/Q _08284_/X _08110_/X _08286_/X _08278_/X vssd1 vssd1 vccd1 vccd1
+ _13930_/D sky130_fd_sc_hd__o221a_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07238_ _07238_/A vssd1 vssd1 vccd1 vccd1 _07238_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07169_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07169_/X sky130_fd_sc_hd__buf_2
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _11648_/A vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__buf_2
XFILLER_133_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput570 _12195_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput581 _13269_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput592 _13279_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13870_ _14107_/CLK _13870_/D vssd1 vssd1 vccd1 vccd1 _13870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12821_ _12517_/X _12820_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12821_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12752_ _09552_/X input339/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ _13648_/Q vssd1 vssd1 vccd1 vccd1 _11703_/Y sky130_fd_sc_hd__inv_2
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12683_ _09589_/X _12682_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13195_/D sky130_fd_sc_hd__mux2_1
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14422_ _14538_/CLK _14422_/D vssd1 vssd1 vccd1 vccd1 _14422_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _13452_/Q vssd1 vssd1 vccd1 vccd1 _11634_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ _14629_/CLK _14353_/D vssd1 vssd1 vccd1 vccd1 _14353_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11565_ _14003_/Q vssd1 vssd1 vccd1 vccd1 _11565_/Y sky130_fd_sc_hd__inv_2
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13304_ _13352_/CLK _13304_/D vssd1 vssd1 vccd1 vccd1 _13304_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10516_ _10510_/Y _10512_/X _10513_/Y _10515_/X vssd1 vssd1 vccd1 vccd1 _10516_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14284_ _14325_/CLK _14284_/D vssd1 vssd1 vccd1 vccd1 _14284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11496_ _14196_/Q vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13235_ _13352_/CLK _13235_/D vssd1 vssd1 vccd1 vccd1 _13267_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _11648_/A vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__buf_4
XFILLER_152_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13166_ _13165_/X _12661_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__mux2_1
X_10378_ _10376_/Y _10248_/X _10377_/Y _10251_/X vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12117_ vssd1 vssd1 vccd1 vccd1 _12117_/HI _12117_/LO sky130_fd_sc_hd__conb_1
XFILLER_170_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13097_ _12627_/X _13096_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12048_ _09781_/A _12043_/X _09893_/A _12044_/X vssd1 vssd1 vccd1 vccd1 _12048_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_22_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13999_ _14110_/CLK _13999_/D vssd1 vssd1 vccd1 vccd1 _13999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06540_ _06540_/A vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__buf_4
XFILLER_74_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_190 input353/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__buf_4
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _09219_/A vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08141_ _13997_/Q _08136_/X _08140_/X _08138_/X _08134_/X vssd1 vssd1 vccd1 vccd1
+ _13997_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08072_ _14026_/Q _08069_/X _07774_/X _08070_/X _08066_/X vssd1 vssd1 vccd1 vccd1
+ _14026_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07023_ _14555_/Q _07014_/X _06725_/X _07017_/X _07018_/X vssd1 vssd1 vccd1 vccd1
+ _14555_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08974_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08974_/X sky130_fd_sc_hd__buf_4
XPHY_7319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput309 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _06495_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07925_ _14106_/Q _07918_/X _07767_/X _07919_/X _07921_/X vssd1 vssd1 vccd1 vccd1
+ _14106_/D sky130_fd_sc_hd__o221a_1
XPHY_6618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07856_ _07856_/A vssd1 vssd1 vccd1 vccd1 _07856_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06807_ _08162_/A vssd1 vssd1 vccd1 vccd1 _06807_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07787_ _14177_/Q _07783_/X _07471_/X _07785_/X _07781_/X vssd1 vssd1 vccd1 vccd1
+ _14177_/D sky130_fd_sc_hd__o221a_1
XFILLER_72_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09526_ _09533_/A _12409_/X vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__and2_1
X_06738_ _07723_/A vssd1 vssd1 vccd1 vccd1 _06738_/X sky130_fd_sc_hd__buf_2
XFILLER_71_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09457_ _09457_/A _12955_/X vssd1 vssd1 vccd1 vccd1 _13287_/D sky130_fd_sc_hd__and2_1
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06669_ _06546_/A _06645_/Y _06544_/Y _08927_/A vssd1 vssd1 vccd1 vccd1 _06669_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _13858_/Q _08344_/A _08268_/X _08346_/A _08406_/X vssd1 vssd1 vccd1 vccd1
+ _13858_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09388_ _09388_/A _13179_/X vssd1 vssd1 vccd1 vccd1 _13343_/D sky130_fd_sc_hd__and2_1
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08339_ _13897_/Q _08274_/A _08268_/X _08276_/A _08336_/X vssd1 vssd1 vccd1 vccd1
+ _13897_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ _14466_/Q vssd1 vssd1 vccd1 vccd1 _11350_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _13658_/Q vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11281_ _13958_/Q vssd1 vssd1 vccd1 vccd1 _11281_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13020_ _12590_/X input354/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13020_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10232_ _14170_/Q vssd1 vssd1 vccd1 vccd1 _10232_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _11830_/A vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10094_ _10094_/A _12481_/X vssd1 vssd1 vccd1 vccd1 _12242_/A sky130_fd_sc_hd__nor2_8
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _14143_/CLK _13922_/D vssd1 vssd1 vccd1 vccd1 _13922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13853_ _14095_/CLK _13853_/D vssd1 vssd1 vccd1 vccd1 _13853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _12513_/X input357/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12804_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13784_ _14121_/CLK _13784_/D vssd1 vssd1 vccd1 vccd1 _13784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10996_ _13672_/Q vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12735_ _09539_/X _12734_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13214_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12666_ _09795_/Y _13343_/Q _12666_/S vssd1 vssd1 vccd1 vccd1 _12666_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _14481_/CLK _14405_/D vssd1 vssd1 vccd1 vccd1 _14405_/Q sky130_fd_sc_hd__dfxtp_1
X_11617_ _11612_/Y _11435_/X _11613_/Y _11437_/X _11616_/X vssd1 vssd1 vccd1 vccd1
+ _11630_/B sky130_fd_sc_hd__o221a_2
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _09917_/X _13314_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12597_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11548_ _11529_/X _11548_/B _11548_/C _11548_/D vssd1 vssd1 vccd1 vccd1 _11549_/D
+ sky130_fd_sc_hd__and4b_1
X_14336_ _14611_/CLK _14336_/D vssd1 vssd1 vccd1 vccd1 _14336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14267_ _14495_/CLK _14267_/D vssd1 vssd1 vccd1 vccd1 _14267_/Q sky130_fd_sc_hd__dfxtp_1
X_11479_ _14118_/Q vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__inv_2
X_13218_ _13350_/CLK _13218_/D vssd1 vssd1 vccd1 vccd1 _13218_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14198_ _14470_/CLK _14198_/D vssd1 vssd1 vccd1 vccd1 _14198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13149_ _12653_/X _13148_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _07710_/A vssd1 vssd1 vccd1 vccd1 _07710_/X sky130_fd_sc_hd__buf_4
XFILLER_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08690_ _13728_/Q _08687_/X _08501_/X _08689_/X _08684_/X vssd1 vssd1 vccd1 vccd1
+ _13728_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07641_ _14244_/Q _07634_/X _07315_/X _07636_/X _07640_/X vssd1 vssd1 vccd1 vccd1
+ _14244_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07572_ _07614_/A vssd1 vssd1 vccd1 vccd1 _07606_/A sky130_fd_sc_hd__buf_4
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09311_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09311_/X sky130_fd_sc_hd__clkbuf_2
X_06523_ _07086_/B vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__inv_2
XFILLER_55_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09242_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ _09173_/A vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__buf_1
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08055_ _14037_/Q _08053_/X _07746_/X _08054_/X _08050_/X vssd1 vssd1 vccd1 vccd1
+ _14037_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07006_ _08989_/B vssd1 vssd1 vccd1 vccd1 _07878_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_162_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput106 la_data_in[45] vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__clkbuf_4
XPHY_7127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput117 la_data_in[55] vssd1 vssd1 vccd1 vccd1 _06553_/A sky130_fd_sc_hd__buf_2
XPHY_7138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput128 la_data_in[65] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput139 la_data_in[75] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__buf_1
XFILLER_44_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _08957_/A vssd1 vssd1 vccd1 vccd1 _08957_/X sky130_fd_sc_hd__buf_4
XPHY_6415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07908_ _14117_/Q _07902_/X _07740_/X _07903_/X _07905_/X vssd1 vssd1 vccd1 vccd1
+ _14117_/D sky130_fd_sc_hd__o221a_1
XPHY_6448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _13618_/Q _08818_/A _08581_/X _08820_/A _08886_/X vssd1 vssd1 vccd1 vccd1
+ _13618_/D sky130_fd_sc_hd__o221a_1
XPHY_6459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10850_ _13871_/Q vssd1 vssd1 vccd1 vccd1 _10850_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _09509_/A _12397_/X vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__and2_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _14376_/Q vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__inv_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12520_ _13364_/Q _10043_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12451_ _12450_/X _06920_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11402_ _13642_/Q vssd1 vssd1 vccd1 vccd1 _11402_/Y sky130_fd_sc_hd__inv_2
X_12382_ _12381_/X _13211_/Q _12645_/S vssd1 vssd1 vccd1 vccd1 _12382_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_90 _08956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14121_ _14121_/CLK _14121_/D vssd1 vssd1 vccd1 vccd1 _14121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ _13562_/Q _11194_/X _13803_/Q _11195_/X vssd1 vssd1 vccd1 vccd1 _11333_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14052_ _14056_/CLK _14052_/D vssd1 vssd1 vccd1 vccd1 _14052_/Q sky130_fd_sc_hd__dfxtp_1
X_11264_ _13918_/Q vssd1 vssd1 vccd1 vccd1 _11264_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13003_ _12580_/X _13002_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13003_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10215_ _14326_/Q vssd1 vssd1 vccd1 vccd1 _10215_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11195_ _11431_/A vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10146_ _10146_/A _12421_/X vssd1 vssd1 vccd1 vccd1 _10146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__or2_2
XFILLER_43_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ _14139_/CLK _13905_/D vssd1 vssd1 vccd1 vccd1 _13905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13836_ _14107_/CLK _13836_/D vssd1 vssd1 vccd1 vccd1 _13836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13767_ _14120_/CLK _13767_/D vssd1 vssd1 vccd1 vccd1 _13767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10979_ _11451_/A vssd1 vssd1 vccd1 vccd1 _10979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12718_ _09569_/X _12717_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13698_ _14169_/CLK _13698_/D vssd1 vssd1 vccd1 vccd1 _13698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _13336_/Q _12648_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14319_ _14637_/CLK _14319_/D vssd1 vssd1 vccd1 vccd1 _14319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09860_ _13308_/Q vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__inv_2
XFILLER_119_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08811_ _13657_/Q _08748_/A _08581_/X _08750_/A _08808_/X vssd1 vssd1 vccd1 vccd1
+ _13657_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09791_ _09791_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__or2_1
XFILLER_140_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08742_ _13695_/Q _08677_/A _08657_/X _08679_/A _08737_/X vssd1 vssd1 vccd1 vccd1
+ _13695_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ _08744_/A _09201_/B _09271_/C _08673_/D vssd1 vssd1 vccd1 vccd1 _10171_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_113_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07624_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07624_/X sky130_fd_sc_hd__buf_2
XPHY_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07555_ _08989_/A vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06506_ _06512_/A vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__inv_2
XFILLER_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07486_ _07542_/A vssd1 vssd1 vccd1 vccd1 _07541_/A sky130_fd_sc_hd__inv_2
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08107_ _14009_/Q _08095_/X _08105_/X _08097_/X _08106_/X vssd1 vssd1 vccd1 vccd1
+ _14009_/D sky130_fd_sc_hd__o221a_1
XFILLER_181_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09087_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08038_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10000_ _13371_/Q _10000_/B vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _09989_/A vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__inv_2
XPHY_6212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11951_ _13693_/Q vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__inv_2
XPHY_6278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _14496_/Q vssd1 vssd1 vccd1 vccd1 _10902_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11882_ _14010_/Q vssd1 vssd1 vccd1 vccd1 _11882_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13621_ _14047_/CLK _13621_/D vssd1 vssd1 vccd1 vccd1 _13621_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10833_ _14143_/Q vssd1 vssd1 vccd1 vccd1 _10833_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10764_ _13947_/Q vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13552_ _14120_/CLK _13552_/D vssd1 vssd1 vccd1 vccd1 _13552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12503_ _12509_/X _06996_/Y _12503_/S vssd1 vssd1 vccd1 vccd1 _12503_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13483_ _14595_/CLK _13483_/D vssd1 vssd1 vccd1 vccd1 _13483_/Q sky130_fd_sc_hd__dfxtp_1
X_10695_ _10686_/Y _10687_/X _10688_/Y _10689_/X _10694_/X vssd1 vssd1 vccd1 vccd1
+ _10755_/A sky130_fd_sc_hd__o221a_1
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12434_ _12509_/X _06902_/Y _12434_/S vssd1 vssd1 vccd1 vccd1 _12434_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12365_ _13200_/Q input97/X _12407_/S vssd1 vssd1 vccd1 vccd1 _12365_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14104_ _14110_/CLK _14104_/D vssd1 vssd1 vccd1 vccd1 _14104_/Q sky130_fd_sc_hd__dfxtp_1
X_11316_ _13679_/Q vssd1 vssd1 vccd1 vccd1 _11316_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ _11507_/Y _14547_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14035_ _14114_/CLK _14035_/D vssd1 vssd1 vccd1 vccd1 _14035_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _11245_/Y _11188_/X _11246_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11247_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11178_ _11414_/A vssd1 vssd1 vccd1 vccd1 _11178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _10137_/A _12445_/X vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13819_ _14095_/CLK _13819_/D vssd1 vssd1 vccd1 vccd1 _13819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07340_ _14392_/Q _07335_/X _07339_/X _07337_/X _07333_/X vssd1 vssd1 vccd1 vccd1
+ _14392_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07271_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07271_/X sky130_fd_sc_hd__buf_2
XFILLER_177_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ _13570_/Q _09004_/X _09009_/X _09006_/X _09000_/X vssd1 vssd1 vccd1 vccd1
+ _13570_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__or2_1
XFILLER_67_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _09843_/A vssd1 vssd1 vccd1 vccd1 _09843_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__or2_1
X_06986_ _06974_/X _12317_/X _06985_/Y _06976_/X vssd1 vssd1 vccd1 vccd1 _06987_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08725_ _13707_/Q _08722_/X _08556_/X _08723_/X _08720_/X vssd1 vssd1 vccd1 vccd1
+ _13707_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08656_ _13742_/Q _08588_/A _08581_/X _08591_/A _08653_/X vssd1 vssd1 vccd1 vccd1
+ _13742_/D sky130_fd_sc_hd__o221a_1
XPHY_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _14261_/Q _07605_/X _07374_/X _07606_/X _07601_/X vssd1 vssd1 vccd1 vccd1
+ _14261_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08587_ _08643_/A vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ _14298_/Q _07532_/X _07379_/X _07533_/X _07536_/X vssd1 vssd1 vccd1 vccd1
+ _14298_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07469_ _07476_/A vssd1 vssd1 vccd1 vccd1 _07469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _13460_/Q _09205_/X _08895_/X _09207_/X _09196_/X vssd1 vssd1 vccd1 vccd1
+ _13460_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _11671_/A vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__buf_2
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09139_ _09173_/A vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12150_ vssd1 vssd1 vccd1 vccd1 _12150_/HI _12150_/LO sky130_fd_sc_hd__conb_1
XFILLER_191_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11101_ _14617_/Q vssd1 vssd1 vccd1 vccd1 _11101_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ vssd1 vssd1 vccd1 vccd1 _12081_/HI _12081_/LO sky130_fd_sc_hd__conb_1
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11032_ _11030_/Y _10987_/X _11031_/Y _10989_/X vssd1 vssd1 vccd1 vccd1 _11032_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12983_ _12570_/X _12982_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12983_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11934_ _11929_/Y _10214_/A _11930_/Y _10217_/A _11933_/X vssd1 vssd1 vccd1 vccd1
+ _11947_/B sky130_fd_sc_hd__o221a_4
XPHY_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11865_ _11846_/X _11865_/B _11865_/C _11865_/D vssd1 vssd1 vccd1 vccd1 _11866_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _14470_/CLK _13604_/D vssd1 vssd1 vccd1 vccd1 _13604_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10816_ _10814_/Y _10714_/X _10815_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _10816_/X
+ sky130_fd_sc_hd__o22a_1
X_11796_ _14125_/Q vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__inv_2
X_14584_ _14621_/CLK _14584_/D vssd1 vssd1 vccd1 vccd1 _14584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13535_ _14130_/CLK _13535_/D vssd1 vssd1 vccd1 vccd1 _13535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _11457_/A vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13466_ _14178_/CLK _13466_/D vssd1 vssd1 vccd1 vccd1 _13466_/Q sky130_fd_sc_hd__dfxtp_1
X_10678_ _13906_/Q vssd1 vssd1 vccd1 vccd1 _10678_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12417_ _13215_/Q _12416_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12417_/X sky130_fd_sc_hd__mux2_1
X_13397_ _14188_/CLK _13397_/D vssd1 vssd1 vccd1 vccd1 _13397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12348_ _13206_/Q _12347_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12348_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12279_ _12071_/Y _13380_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _14121_/CLK _14018_/D vssd1 vssd1 vccd1 vccd1 _14018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06840_ _08981_/A vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__buf_4
XFILLER_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06771_ _08137_/A vssd1 vssd1 vccd1 vccd1 _06771_/X sky130_fd_sc_hd__buf_2
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08510_ _08914_/A vssd1 vssd1 vccd1 vccd1 _08510_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ _13269_/Q _09486_/X _12264_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _13269_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08441_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08372_ _08389_/A vssd1 vssd1 vccd1 vccd1 _08372_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07323_ _07719_/A vssd1 vssd1 vccd1 vccd1 _07323_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07254_ _07262_/A vssd1 vssd1 vccd1 vccd1 _07254_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07185_ _07209_/A vssd1 vssd1 vccd1 vccd1 _07185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09826_ _13338_/Q _09824_/Y _09789_/B vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09757_ _13331_/Q vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__inv_2
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06969_ _06972_/A _06969_/B vssd1 vssd1 vccd1 vccd1 _14570_/D sky130_fd_sc_hd__nor2_1
XFILLER_189_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08708_ _13718_/Q _08706_/X _08527_/X _08707_/X _08704_/X vssd1 vssd1 vccd1 vccd1
+ _13718_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09688_ _14573_/Q _06964_/Y _06957_/Y _14571_/Q vssd1 vssd1 vccd1 vccd1 _09688_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _13753_/Q _08635_/X _08556_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _13753_/D sky130_fd_sc_hd__o221a_1
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11650_ _11650_/A vssd1 vssd1 vccd1 vccd1 _11650_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _10596_/Y _10506_/X _10597_/Y _10509_/X _10600_/X vssd1 vssd1 vccd1 vccd1
+ _10602_/D sky130_fd_sc_hd__o221a_1
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _11579_/Y _11449_/X _11580_/Y _11451_/X vssd1 vssd1 vccd1 vccd1 _11581_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _13825_/Q vssd1 vssd1 vccd1 vccd1 _10532_/Y sky130_fd_sc_hd__inv_2
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _13352_/CLK _13320_/D vssd1 vssd1 vccd1 vccd1 _13320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10463_ _13505_/Q vssd1 vssd1 vccd1 vccd1 _10463_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13251_ _13372_/CLK _13251_/D vssd1 vssd1 vccd1 vccd1 _13283_/Q sky130_fd_sc_hd__dfxtp_4
X_12202_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _14589_/Q _14590_/Q _14587_/Q _14588_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13182_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10394_ _13823_/Q vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12133_ vssd1 vssd1 vccd1 vccd1 _12133_/HI _12133_/LO sky130_fd_sc_hd__conb_1
XFILLER_135_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12064_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11015_ _13207_/Q _11013_/X _14030_/Q _10957_/X _11014_/X vssd1 vssd1 vccd1 vccd1
+ _11015_/X sky130_fd_sc_hd__a221o_4
XFILLER_113_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12966_ _12965_/X _12562_/X _12974_/S vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11917_ _13777_/Q vssd1 vssd1 vccd1 vccd1 _11917_/Y sky130_fd_sc_hd__inv_2
XPHY_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12535_/X _12896_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12897_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14636_ _14637_/CLK _14636_/D vssd1 vssd1 vccd1 vccd1 _14636_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _14360_/Q vssd1 vssd1 vccd1 vccd1 _11848_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ _14573_/CLK _14567_/D vssd1 vssd1 vccd1 vccd1 _14567_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11779_ _11777_/Y _11693_/X _11778_/Y _11695_/X vssd1 vssd1 vccd1 vccd1 _11779_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13518_ _14110_/CLK _13518_/D vssd1 vssd1 vccd1 vccd1 _13518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14498_ _14621_/CLK _14498_/D vssd1 vssd1 vccd1 vccd1 _14498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13449_ _14183_/CLK _13449_/D vssd1 vssd1 vccd1 vccd1 _13449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ _09132_/A _10204_/A vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__or2_2
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07941_ _14099_/Q _07934_/X _07867_/X _07935_/X _07940_/X vssd1 vssd1 vccd1 vccd1
+ _14099_/D sky130_fd_sc_hd__o221a_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07872_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07872_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_211_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09611_ _14593_/Q _06964_/Y _06881_/Y _14571_/Q vssd1 vssd1 vccd1 vccd1 _09611_/X
+ sky130_fd_sc_hd__a22o_1
X_06823_ _06823_/A vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06754_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06754_/X sky130_fd_sc_hd__clkbuf_2
X_09542_ _09530_/X _09541_/X _13277_/Q _09531_/X vssd1 vssd1 vccd1 vccd1 _13245_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09473_ _09480_/A vssd1 vssd1 vccd1 vccd1 _09473_/X sky130_fd_sc_hd__clkbuf_2
X_06685_ _06562_/A _06684_/X _06562_/A _06684_/X vssd1 vssd1 vccd1 vccd1 _06685_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08424_ _08468_/A vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08355_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07306_ _07387_/A vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08286_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07237_ _07290_/A vssd1 vssd1 vccd1 vccd1 _07238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07168_ _14480_/Q _07164_/X _06714_/X _07166_/X _07153_/X vssd1 vssd1 vccd1 vccd1
+ _14480_/D sky130_fd_sc_hd__o221a_1
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07099_ _14517_/Q _07092_/X _06722_/X _07094_/X _07096_/X vssd1 vssd1 vccd1 vccd1
+ _14517_/D sky130_fd_sc_hd__o221a_1
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput560 _12186_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput571 _12232_/X vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput582 _13270_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput593 _13280_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09809_ _09812_/B vssd1 vssd1 vccd1 vccd1 _09809_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12820_ _12517_/X input341/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12751_ _09550_/X _12750_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13210_/D sky130_fd_sc_hd__mux2_1
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _13687_/Q vssd1 vssd1 vccd1 vccd1 _11702_/Y sky130_fd_sc_hd__inv_2
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _09589_/X _12681_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12682_/X sky130_fd_sc_hd__mux2_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14459_/CLK _14421_/D vssd1 vssd1 vccd1 vccd1 _14421_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A vssd1 vssd1 vccd1 vccd1 _11633_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14352_ _14629_/CLK _14352_/D vssd1 vssd1 vccd1 vccd1 _14352_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11564_ _11562_/Y _11419_/X _11563_/Y _11421_/X vssd1 vssd1 vccd1 vccd1 _11564_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13303_ _13352_/CLK _13303_/D vssd1 vssd1 vccd1 vccd1 _13303_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10515_ _11461_/A vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14283_ _14325_/CLK _14283_/D vssd1 vssd1 vccd1 vccd1 _14283_/Q sky130_fd_sc_hd__dfxtp_1
X_11495_ _13604_/Q vssd1 vssd1 vccd1 vccd1 _11495_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10446_ _13746_/Q vssd1 vssd1 vccd1 vccd1 _10446_/Y sky130_fd_sc_hd__inv_2
X_13234_ _13352_/CLK _13234_/D vssd1 vssd1 vccd1 vccd1 _13266_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10377_ _14446_/Q vssd1 vssd1 vccd1 vccd1 _10377_/Y sky130_fd_sc_hd__inv_2
X_13165_ _12661_/X _13164_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12116_ vssd1 vssd1 vccd1 vccd1 _12116_/HI _12116_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13096_ _12627_/X input333/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _09780_/A _12043_/X _09892_/A _12044_/X vssd1 vssd1 vccd1 vccd1 _12047_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_26_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13998_ _14120_/CLK _13998_/D vssd1 vssd1 vccd1 vccd1 _13998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12949_ _12555_/X _12948_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_180 input334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_191 input355/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ _14621_/CLK _14619_/D vssd1 vssd1 vccd1 vccd1 _14619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _08140_/A vssd1 vssd1 vccd1 vccd1 _08140_/X sky130_fd_sc_hd__buf_4
XFILLER_159_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08071_ _14027_/Q _08069_/X _07771_/X _08070_/X _08066_/X vssd1 vssd1 vccd1 vccd1
+ _14027_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07022_ _14556_/Q _07014_/X _06722_/X _07017_/X _07018_/X vssd1 vssd1 vccd1 vccd1
+ _14556_/D sky130_fd_sc_hd__o221a_1
XFILLER_122_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08973_ _13585_/Q _08969_/X _08648_/X _08971_/X _08963_/X vssd1 vssd1 vccd1 vccd1
+ _13585_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07924_ _14107_/Q _07918_/X _07852_/X _07919_/X _07921_/X vssd1 vssd1 vccd1 vccd1
+ _14107_/D sky130_fd_sc_hd__o221a_1
XPHY_6608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07855_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06806_ _08957_/A vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07786_ _14178_/Q _07783_/X _07784_/X _07785_/X _07781_/X vssd1 vssd1 vccd1 vccd1
+ _14178_/D sky130_fd_sc_hd__o221a_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _09514_/X _09524_/X _13283_/Q _09517_/X vssd1 vssd1 vccd1 vccd1 _13251_/D
+ sky130_fd_sc_hd__o22a_1
X_06737_ _08837_/A vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06668_ _06668_/A vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__buf_2
X_09456_ _09456_/A _12951_/X vssd1 vssd1 vccd1 vccd1 _13288_/D sky130_fd_sc_hd__and2_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _13859_/Q _08344_/A _08190_/X _08346_/A _08406_/X vssd1 vssd1 vccd1 vccd1
+ _13859_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06599_ _06540_/A _06598_/A _06538_/Y _06598_/Y vssd1 vssd1 vccd1 vccd1 _06599_/X
+ sky130_fd_sc_hd__a22o_1
X_09387_ _09388_/A _13175_/X vssd1 vssd1 vccd1 vccd1 _13344_/D sky130_fd_sc_hd__and2_1
XFILLER_71_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08338_ _13898_/Q _08274_/A _08190_/X _08276_/A _08336_/X vssd1 vssd1 vccd1 vccd1
+ _13898_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08269_ _13936_/Q _08198_/A _08268_/X _08201_/A _08264_/X vssd1 vssd1 vccd1 vccd1
+ _13936_/D sky130_fd_sc_hd__o221a_1
XFILLER_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10300_ _13424_/Q vssd1 vssd1 vccd1 vccd1 _10300_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ _14231_/Q _11170_/X _14426_/Q _11171_/X _11279_/X vssd1 vssd1 vccd1 vccd1
+ _11313_/B sky130_fd_sc_hd__a221oi_2
XFILLER_88_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ _10231_/A vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10162_/A vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__inv_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput390 _12198_/X vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10093_ _10099_/A _10134_/A vssd1 vssd1 vccd1 vccd1 _12479_/S sky130_fd_sc_hd__or2_1
XFILLER_47_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13921_ _14143_/CLK _13921_/D vssd1 vssd1 vccd1 vccd1 _13921_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13852_ _14094_/CLK _13852_/D vssd1 vssd1 vccd1 vccd1 _13852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12803_ _12512_/X _12802_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13783_ _14123_/CLK _13783_/D vssd1 vssd1 vccd1 vccd1 _13783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10995_ _13438_/Q vssd1 vssd1 vccd1 vccd1 _10995_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ _09539_/X _12733_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12734_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _13344_/Q _12664_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12665_/X sky130_fd_sc_hd__mux2_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14481_/CLK _14404_/D vssd1 vssd1 vccd1 vccd1 _14404_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _11614_/Y _11439_/X _11615_/Y _11441_/X vssd1 vssd1 vccd1 vccd1 _11616_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12596_ _13315_/Q _12595_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12596_/X sky130_fd_sc_hd__mux2_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14335_ _14611_/CLK _14335_/D vssd1 vssd1 vccd1 vccd1 _14335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11547_ _11542_/Y _11455_/X _11543_/Y _11457_/X _11546_/X vssd1 vssd1 vccd1 vccd1
+ _11548_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14266_ _14305_/CLK _14266_/D vssd1 vssd1 vccd1 vccd1 _14266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11478_ _13845_/Q vssd1 vssd1 vccd1 vccd1 _11478_/Y sky130_fd_sc_hd__inv_2
X_13217_ _14459_/CLK _13217_/D vssd1 vssd1 vccd1 vccd1 _13217_/Q sky130_fd_sc_hd__dfxtp_4
X_10429_ _13661_/Q vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _14470_/CLK _14197_/D vssd1 vssd1 vccd1 vccd1 _14197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13148_ _12653_/X input354/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13079_ _12618_/X _13078_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07640_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07640_/X sky130_fd_sc_hd__buf_2
XFILLER_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07571_ _07605_/A vssd1 vssd1 vccd1 vccd1 _07571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06522_ _08482_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09310_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09241_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09172_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _08123_/A vssd1 vssd1 vccd1 vccd1 _08123_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07005_ _07803_/A vssd1 vssd1 vccd1 vccd1 _07484_/A sky130_fd_sc_hd__buf_1
XFILLER_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 la_data_in[46] vssd1 vssd1 vccd1 vccd1 _06614_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 la_data_in[56] vssd1 vssd1 vccd1 vccd1 _06595_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08956_ _08956_/A vssd1 vssd1 vccd1 vccd1 _08956_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput129 la_data_in[66] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__buf_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07907_ _14118_/Q _07902_/X _07738_/X _07903_/X _07905_/X vssd1 vssd1 vccd1 vccd1
+ _14118_/D sky130_fd_sc_hd__o221a_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _13619_/Q _08818_/A _08579_/X _08820_/A _08886_/X vssd1 vssd1 vccd1 vccd1
+ _13619_/D sky130_fd_sc_hd__o221a_1
XPHY_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _07856_/A vssd1 vssd1 vccd1 vccd1 _07838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07769_ _14184_/Q _07758_/X _07767_/X _07760_/X _07768_/X vssd1 vssd1 vccd1 vccd1
+ _14184_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ _13255_/Q _09479_/A _12250_/X _09480_/A vssd1 vssd1 vccd1 vccd1 _13255_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _14610_/Q vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09445_/A vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__clkbuf_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12450_ _12449_/X _06920_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11401_ _11401_/A vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12381_ _13211_/Q _12380_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12381_/X sky130_fd_sc_hd__mux2_1
XANTENNA_80 _08183_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_91 _08958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14120_ _14120_/CLK _14120_/D vssd1 vssd1 vccd1 vccd1 _14120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11332_ _11322_/Y _11176_/X _11325_/X _11328_/X _11331_/X vssd1 vssd1 vccd1 vccd1
+ _11354_/C sky130_fd_sc_hd__o2111a_4
XFILLER_193_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14051_ _14056_/CLK _14051_/D vssd1 vssd1 vccd1 vccd1 _14051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11263_ _11258_/Y _11209_/X _11259_/Y _11211_/X _11262_/X vssd1 vssd1 vccd1 vccd1
+ _11270_/C sky130_fd_sc_hd__o221a_1
XFILLER_175_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _13001_/X _12580_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10214_ _10214_/A vssd1 vssd1 vccd1 vccd1 _10214_/X sky130_fd_sc_hd__clkbuf_2
X_11194_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _12419_/S sky130_fd_sc_hd__or2_1
XFILLER_121_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10076_ _10076_/A _12496_/X vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__nor2_8
XFILLER_43_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _14139_/CLK _13904_/D vssd1 vssd1 vccd1 vccd1 _13904_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13835_ _14107_/CLK _13835_/D vssd1 vssd1 vccd1 vccd1 _13835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13766_ _14120_/CLK _13766_/D vssd1 vssd1 vccd1 vccd1 _13766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10978_ _14263_/Q vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12717_ _09569_/X _12716_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13697_ _14173_/CLK _13697_/D vssd1 vssd1 vccd1 vccd1 _13697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _09823_/X _13336_/Q _12650_/S vssd1 vssd1 vccd1 vccd1 _12648_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _09938_/Y _13307_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14318_ _14481_/CLK _14318_/D vssd1 vssd1 vccd1 vccd1 _14318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14249_ _14325_/CLK _14249_/D vssd1 vssd1 vccd1 vccd1 _14249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08810_ _13658_/Q _08748_/A _08579_/X _08750_/A _08808_/X vssd1 vssd1 vccd1 vccd1
+ _13658_/D sky130_fd_sc_hd__o221a_1
X_09790_ _09790_/A _09827_/A vssd1 vssd1 vccd1 vccd1 _09791_/B sky130_fd_sc_hd__or2_2
XFILLER_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08741_ _13696_/Q _08677_/A _08581_/X _08679_/A _08737_/X vssd1 vssd1 vccd1 vccd1
+ _13696_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08672_ _13734_/Q _08662_/A _08505_/X _08663_/A _08671_/X vssd1 vssd1 vccd1 vccd1
+ _13734_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07623_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07554_ _07803_/A vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__inv_2
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06505_ _06507_/A _06507_/B _06507_/C _06508_/A vssd1 vssd1 vccd1 vccd1 _06505_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_165_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07485_ _07558_/A _11679_/A vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__or2_2
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09224_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09155_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08106_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08106_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09086_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ _08079_/A vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__buf_2
XFILLER_102_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _13365_/Q _09988_/B vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08939_ _13599_/Q _08929_/X _08935_/X _08931_/X _08938_/X vssd1 vssd1 vccd1 vccd1
+ _13599_/D sky130_fd_sc_hd__o221a_1
XPHY_6235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11950_ _13459_/Q vssd1 vssd1 vccd1 vccd1 _11950_/Y sky130_fd_sc_hd__inv_2
XPHY_6268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater690 _12647_/S vssd1 vssd1 vccd1 vccd1 _12645_/S sky130_fd_sc_hd__buf_8
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10901_ _13205_/Q _10775_/X _14028_/Q _10719_/X _10900_/X vssd1 vssd1 vccd1 vccd1
+ _10901_/X sky130_fd_sc_hd__a221o_2
XPHY_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11881_ _11879_/Y _10188_/A _11880_/Y _10191_/A vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13620_ _14047_/CLK _13620_/D vssd1 vssd1 vccd1 vccd1 _13620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10832_ _13909_/Q vssd1 vssd1 vccd1 vccd1 _10832_/Y sky130_fd_sc_hd__inv_2
XPHY_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13551_ _14120_/CLK _13551_/D vssd1 vssd1 vccd1 vccd1 _13551_/Q sky130_fd_sc_hd__dfxtp_1
X_10763_ _14220_/Q _10696_/X _14415_/Q _10697_/X _10762_/X vssd1 vssd1 vccd1 vccd1
+ _10797_/B sky130_fd_sc_hd__a221oi_2
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12502_ _12501_/X _06989_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__mux2_2
XFILLER_185_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13482_ _14595_/CLK _13482_/D vssd1 vssd1 vccd1 vccd1 _13482_/Q sky130_fd_sc_hd__dfxtp_1
X_10694_ _10690_/Y _10691_/X _10692_/Y _10693_/X vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ _12432_/X _06897_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12433_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ _12363_/X _13201_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12364_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14103_ _14110_/CLK _14103_/D vssd1 vssd1 vccd1 vccd1 _14103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11315_ _13445_/Q vssd1 vssd1 vccd1 vccd1 _11315_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ _11549_/Y _14548_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__mux2_2
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14034_ _14114_/CLK _14034_/D vssd1 vssd1 vccd1 vccd1 _14034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11246_ _13521_/Q vssd1 vssd1 vccd1 vccd1 _11246_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11177_ _13761_/Q vssd1 vssd1 vccd1 vccd1 _11177_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10128_ _10128_/A vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10059_ _10081_/A vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__buf_1
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ _14130_/CLK _13818_/D vssd1 vssd1 vccd1 vccd1 _13818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13749_ _14121_/CLK _13749_/D vssd1 vssd1 vccd1 vccd1 _13749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07270_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__buf_4
XFILLER_182_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09911_ _13313_/Q vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__inv_2
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09842_ _13332_/Q _09840_/Y _09783_/B vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09773_ _09773_/A _09850_/A vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__or2_2
XFILLER_26_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06985_ _14565_/Q vssd1 vssd1 vccd1 vccd1 _06985_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _13708_/Q _08722_/X _08553_/X _08723_/X _08720_/X vssd1 vssd1 vccd1 vccd1
+ _13708_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08655_ _13743_/Q _08588_/A _08579_/X _08591_/A _08653_/X vssd1 vssd1 vccd1 vccd1
+ _13743_/D sky130_fd_sc_hd__o221a_1
XPHY_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07606_ _07606_/A vssd1 vssd1 vccd1 vccd1 _07606_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08586_ _08644_/A vssd1 vssd1 vccd1 vccd1 _08643_/A sky130_fd_sc_hd__inv_2
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07537_ _14299_/Q _07532_/X _07377_/X _07533_/X _07536_/X vssd1 vssd1 vccd1 vccd1
+ _14299_/D sky130_fd_sc_hd__o221a_1
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07468_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07468_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09207_ _09207_/A vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07399_ _08186_/A vssd1 vssd1 vccd1 vccd1 _07399_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ _09138_/A vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__buf_6
XFILLER_202_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09069_/A vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11100_ _14344_/Q vssd1 vssd1 vccd1 vccd1 _11100_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ vssd1 vssd1 vccd1 vccd1 _12080_/HI _12080_/LO sky130_fd_sc_hd__conb_1
XFILLER_172_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11031_ _14459_/Q vssd1 vssd1 vccd1 vccd1 _11031_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12982_ _12981_/X _12570_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _12982_/X sky130_fd_sc_hd__mux2_1
XPHY_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11931_/Y _10220_/A _11932_/Y _10223_/A vssd1 vssd1 vccd1 vccd1 _11933_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _11859_/Y _11689_/X _11860_/Y _11691_/X _11863_/X vssd1 vssd1 vccd1 vccd1
+ _11865_/D sky130_fd_sc_hd__o221a_1
XPHY_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _14470_/CLK _13603_/D vssd1 vssd1 vccd1 vccd1 _13603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _13512_/Q vssd1 vssd1 vccd1 vccd1 _10815_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14583_ _14621_/CLK _14583_/D vssd1 vssd1 vccd1 vccd1 _14583_/Q sky130_fd_sc_hd__dfxtp_2
X_11795_ _13852_/Q vssd1 vssd1 vccd1 vccd1 _11795_/Y sky130_fd_sc_hd__inv_2
XPHY_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13534_ _14130_/CLK _13534_/D vssd1 vssd1 vccd1 vccd1 _13534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _14141_/Q vssd1 vssd1 vccd1 vccd1 _10746_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _14178_/CLK _13465_/D vssd1 vssd1 vccd1 vccd1 _13465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10677_ _10672_/Y _10492_/X _10673_/Y _10495_/X _10676_/X vssd1 vssd1 vccd1 vccd1
+ _10684_/C sky130_fd_sc_hd__o221a_1
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12416_ _13215_/Q _06668_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12416_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _14183_/CLK _13396_/D vssd1 vssd1 vccd1 vccd1 _13396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12347_ _13206_/Q _06703_/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _12070_/Y _13379_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12278_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14017_ _14047_/CLK _14017_/D vssd1 vssd1 vccd1 vccd1 _14017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11229_ _11229_/A _11229_/B _11229_/C _11229_/D vssd1 vssd1 vccd1 vccd1 _11229_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06770_ _08930_/A vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__buf_4
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput290 la_oenb[96] vssd1 vssd1 vccd1 vccd1 input290/X sky130_fd_sc_hd__buf_1
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08440_ _13845_/Q _08436_/X _08128_/X _08437_/X _08433_/X vssd1 vssd1 vccd1 vccd1
+ _13845_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08371_ _08388_/A vssd1 vssd1 vccd1 vccd1 _08371_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07322_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07253_ _14435_/Q _07248_/X _07031_/X _07250_/X _07244_/X vssd1 vssd1 vccd1 vccd1
+ _14435_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07184_ _14472_/Q _07174_/X _06748_/X _07176_/X _07181_/X vssd1 vssd1 vccd1 vccd1
+ _14472_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _09787_/A _09787_/B _09824_/Y vssd1 vssd1 vccd1 vccd1 _09825_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09756_ _13332_/Q vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__inv_2
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06968_ _06956_/X _12312_/X _06967_/Y _06958_/X vssd1 vssd1 vccd1 vccd1 _06969_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08707_ _08723_/A vssd1 vssd1 vccd1 vccd1 _08707_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09687_ _06865_/X _09640_/A _14597_/Q _09640_/Y vssd1 vssd1 vccd1 vccd1 _09687_/X
+ sky130_fd_sc_hd__o22a_1
X_06899_ _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _14589_/D sky130_fd_sc_hd__nor2_1
XFILLER_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _13754_/Q _08635_/X _08553_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _13754_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08569_ _13787_/Q _08565_/X _08259_/X _08567_/X _08563_/X vssd1 vssd1 vccd1 vccd1
+ _13787_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ _10598_/Y _10512_/X _10599_/Y _10515_/X vssd1 vssd1 vccd1 vccd1 _10600_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _14276_/Q vssd1 vssd1 vccd1 vccd1 _11580_/Y sky130_fd_sc_hd__inv_2
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10531_ _10529_/Y _10448_/X _10530_/Y _10451_/X vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13250_ _13372_/CLK _13250_/D vssd1 vssd1 vccd1 vccd1 _13282_/Q sky130_fd_sc_hd__dfxtp_4
X_10462_ _11424_/A vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12201_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13181_ _14577_/Q _14578_/Q _14575_/Q _14576_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13181_/X sky130_fd_sc_hd__mux4_2
XFILLER_174_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10393_ _10391_/Y _10181_/X _10392_/Y _10184_/X vssd1 vssd1 vccd1 vccd1 _10393_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12132_ vssd1 vssd1 vccd1 vccd1 _12132_/HI _12132_/LO sky130_fd_sc_hd__conb_1
XFILLER_174_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _09792_/A _12057_/X _09904_/A _12058_/X vssd1 vssd1 vccd1 vccd1 _12063_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11014_ _13555_/Q _10958_/X _13796_/Q _10959_/X vssd1 vssd1 vccd1 vccd1 _11014_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12965_ _12562_/X _12964_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12965_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11916_ _13972_/Q vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__inv_2
XPHY_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12535_/X input353/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14637_/CLK _14635_/D vssd1 vssd1 vccd1 vccd1 _14635_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ _14516_/Q vssd1 vssd1 vccd1 vccd1 _11847_/Y sky130_fd_sc_hd__inv_2
XPHY_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _14573_/CLK _14566_/D vssd1 vssd1 vccd1 vccd1 _14566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11778_ _14475_/Q vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13517_ _13996_/CLK _13517_/D vssd1 vssd1 vccd1 vccd1 _13517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10729_ _11439_/A vssd1 vssd1 vccd1 vccd1 _10729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14497_ _14621_/CLK _14497_/D vssd1 vssd1 vccd1 vccd1 _14497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13448_ _14183_/CLK _13448_/D vssd1 vssd1 vccd1 vccd1 _13448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13379_ _14538_/CLK _13379_/D vssd1 vssd1 vccd1 vccd1 _13379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07940_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07871_ _14135_/Q _07863_/X _07792_/X _07864_/X _07865_/X vssd1 vssd1 vccd1 vccd1
+ _14135_/D sky130_fd_sc_hd__o221a_1
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09610_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06822_ _14608_/Q _06805_/X _06820_/X _06811_/X _06821_/X vssd1 vssd1 vccd1 vccd1
+ _14608_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09541_ _09547_/A _12376_/X vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__and2_1
XFILLER_168_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06753_ _08123_/A vssd1 vssd1 vccd1 vccd1 _06753_/X sky130_fd_sc_hd__buf_2
XFILLER_97_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09472_ _09479_/A vssd1 vssd1 vccd1 vccd1 _09472_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06684_ _06656_/Y _08960_/A _06657_/A _06559_/Y vssd1 vssd1 vccd1 vccd1 _06684_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08423_ _13853_/Q _08415_/X _08105_/X _08417_/X _08421_/X vssd1 vssd1 vccd1 vccd1
+ _13853_/D sky130_fd_sc_hd__o221a_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08354_ _08388_/A vssd1 vssd1 vccd1 vccd1 _08354_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07305_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__inv_2
XFILLER_123_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08285_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_203_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07236_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07290_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07167_ _14481_/Q _07164_/X _07015_/X _07166_/X _07153_/X vssd1 vssd1 vccd1 vccd1
+ _14481_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07098_ _14518_/Q _07092_/X _06719_/X _07094_/X _07096_/X vssd1 vssd1 vccd1 vccd1
+ _14518_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput550 _12177_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput561 _12187_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__clkbuf_2
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput572 _12233_/X vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput583 _13271_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput594 _13281_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__or2_2
XFILLER_210_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _10112_/A _10081_/A vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__or2_1
XFILLER_95_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12750_ _09550_/X _12749_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12750_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _13453_/Q vssd1 vssd1 vccd1 vccd1 _11701_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12681_ _09589_/X _12680_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12681_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14420_ _14459_/CLK _14420_/D vssd1 vssd1 vccd1 vccd1 _14420_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _14083_/Q vssd1 vssd1 vccd1 vccd1 _11632_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14351_ _14629_/CLK _14351_/D vssd1 vssd1 vccd1 vccd1 _14351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11563_ _14120_/Q vssd1 vssd1 vccd1 vccd1 _11563_/Y sky130_fd_sc_hd__inv_2
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _13352_/CLK _13302_/D vssd1 vssd1 vccd1 vccd1 _13302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _11695_/A vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__buf_4
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _14325_/CLK _14282_/D vssd1 vssd1 vccd1 vccd1 _14282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _14313_/Q vssd1 vssd1 vccd1 vccd1 _11494_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _13352_/CLK _13233_/D vssd1 vssd1 vccd1 vccd1 _13265_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10445_ _11412_/A vssd1 vssd1 vccd1 vccd1 _10445_/X sky130_fd_sc_hd__buf_2
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13164_ _12661_/X input349/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__mux2_1
X_10376_ _13464_/Q vssd1 vssd1 vccd1 vccd1 _10376_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12115_ vssd1 vssd1 vccd1 vccd1 _12115_/HI _12115_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13095_ _12625_/X _13094_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13095_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12046_ _09779_/A _12043_/X _09891_/A _12044_/X vssd1 vssd1 vccd1 vccd1 _12046_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13997_ _14120_/CLK _13997_/D vssd1 vssd1 vccd1 vccd1 _13997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12948_ _12555_/X input341/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _12530_/X _12878_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__mux2_1
XANTENNA_170 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_181 input334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_192 input355/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14618_ _14627_/CLK _14618_/D vssd1 vssd1 vccd1 vccd1 _14618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14549_ _14611_/CLK _14549_/D vssd1 vssd1 vccd1 vccd1 _14549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08070_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08070_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07021_ _14557_/Q _07014_/X _06719_/X _07017_/X _07018_/X vssd1 vssd1 vccd1 vccd1
+ _14557_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08972_ _13586_/Q _08969_/X _08970_/X _08971_/X _08963_/X vssd1 vssd1 vccd1 vccd1
+ _13586_/D sky130_fd_sc_hd__o221a_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07923_ _14108_/Q _07918_/X _07764_/X _07919_/X _07921_/X vssd1 vssd1 vccd1 vccd1
+ _14108_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07854_ _14145_/Q _07845_/X _07767_/X _07846_/X _07848_/X vssd1 vssd1 vccd1 vccd1
+ _14145_/D sky130_fd_sc_hd__o221a_1
XPHY_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06805_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06805_/X sky130_fd_sc_hd__clkbuf_2
X_07785_ _07785_/A vssd1 vssd1 vccd1 vccd1 _07785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09524_ _09533_/A _12406_/X vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__and2_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06736_ _14632_/Q _06733_/X _06735_/X _06726_/X _06730_/X vssd1 vssd1 vccd1 vccd1
+ _14632_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09456_/A _12947_/X vssd1 vssd1 vccd1 vccd1 _13289_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06667_ _06664_/X _06666_/X _06664_/X _06666_/X vssd1 vssd1 vccd1 vccd1 _06667_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _08421_/A vssd1 vssd1 vccd1 vccd1 _08406_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _09388_/A _13171_/X vssd1 vssd1 vccd1 vccd1 _13345_/D sky130_fd_sc_hd__and2_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06598_ _06598_/A vssd1 vssd1 vccd1 vccd1 _06598_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08337_ _13899_/Q _08274_/A _08188_/X _08276_/A _08336_/X vssd1 vssd1 vccd1 vccd1
+ _13899_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08268_ _08268_/A vssd1 vssd1 vccd1 vccd1 _08268_/X sky130_fd_sc_hd__buf_4
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _14451_/Q _07217_/X _06825_/X _07218_/X _07213_/X vssd1 vssd1 vccd1 vccd1
+ _14451_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08199_ _08895_/A vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10230_ _11681_/A vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10148_/Y _10150_/X _10151_/Y _10153_/X _10160_/X vssd1 vssd1 vccd1 vccd1
+ _10255_/A sky130_fd_sc_hd__o221a_2
XFILLER_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _12216_/X vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_175_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput391 _12226_/X vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10102_/B _10132_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__or2_1
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _14146_/CLK _13920_/D vssd1 vssd1 vccd1 vccd1 _13920_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13851_ _14094_/CLK _13851_/D vssd1 vssd1 vccd1 vccd1 _13851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12802_ _12512_/X _12801_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13782_ _14123_/CLK _13782_/D vssd1 vssd1 vccd1 vccd1 _13782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _14069_/Q vssd1 vssd1 vccd1 vccd1 _10994_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12733_ _09539_/X _12732_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12733_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12664_ _09799_/X _13344_/Q _12666_/S vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14403_ _14633_/CLK _14403_/D vssd1 vssd1 vccd1 vccd1 _14403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ _14394_/Q vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__inv_2
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _09921_/Y _13315_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__mux2_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _14527_/CLK _14334_/D vssd1 vssd1 vccd1 vccd1 _14334_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _11544_/Y _11459_/X _11545_/Y _11461_/X vssd1 vssd1 vccd1 vccd1 _11546_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14265_ _14305_/CLK _14265_/D vssd1 vssd1 vccd1 vccd1 _14265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11477_ _11475_/Y _11414_/X _11476_/Y _11416_/X vssd1 vssd1 vccd1 vccd1 _11477_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13216_ _13350_/CLK _13216_/D vssd1 vssd1 vccd1 vccd1 _13216_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10428_ _11399_/A vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14196_ _14529_/CLK _14196_/D vssd1 vssd1 vccd1 vccd1 _14196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _12651_/X _13146_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10359_ _10349_/Y _10178_/X _10352_/X _10355_/X _10358_/X vssd1 vssd1 vccd1 vccd1
+ _10381_/C sky130_fd_sc_hd__o2111a_4
XFILLER_151_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ _13077_/X _12618_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12029_ _12010_/X _12029_/B _12029_/C _12029_/D vssd1 vssd1 vccd1 vccd1 _12030_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_6_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07570_ _07613_/A vssd1 vssd1 vccd1 vccd1 _07605_/A sky130_fd_sc_hd__buf_4
XFILLER_4_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06521_ _08989_/B vssd1 vssd1 vccd1 vccd1 _08482_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09240_ _13441_/Q _09233_/X _08942_/X _09234_/X _09236_/X vssd1 vssd1 vccd1 vccd1
+ _13441_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09171_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08122_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08053_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08053_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ _07004_/A _07004_/B vssd1 vssd1 vccd1 vccd1 _14560_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 la_data_in[47] vssd1 vssd1 vccd1 vccd1 _06554_/A sky130_fd_sc_hd__clkbuf_2
X_08955_ _13592_/Q _08944_/X _08954_/X _08946_/X _08951_/X vssd1 vssd1 vccd1 vccd1
+ _13592_/D sky130_fd_sc_hd__o221a_1
XPHY_7129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput119 la_data_in[57] vssd1 vssd1 vccd1 vccd1 _06611_/A sky130_fd_sc_hd__buf_2
XFILLER_29_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _14119_/Q _07902_/X _07736_/X _07903_/X _07905_/X vssd1 vssd1 vccd1 vccd1
+ _14119_/D sky130_fd_sc_hd__o221a_1
XPHY_6428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _08923_/A vssd1 vssd1 vccd1 vccd1 _08886_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07837_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07837_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07768_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09507_ _13256_/Q _09479_/A _12251_/X _09480_/A vssd1 vssd1 vccd1 vccd1 _13256_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06719_ _07710_/A vssd1 vssd1 vccd1 vccd1 _06719_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07699_ _14209_/Q _07634_/A _07480_/X _07636_/A _07698_/X vssd1 vssd1 vccd1 vccd1
+ _14209_/D sky130_fd_sc_hd__o221a_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _13019_/X vssd1 vssd1 vccd1 vccd1 _13303_/D sky130_fd_sc_hd__and2_1
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09369_ _09370_/A _12859_/X vssd1 vssd1 vccd1 vccd1 _13359_/D sky130_fd_sc_hd__and2_1
XFILLER_51_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ _13681_/Q vssd1 vssd1 vccd1 vccd1 _11400_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12380_ _13211_/Q _06554_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_70 _08155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_81 _08264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_92 _08935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11329_/Y _11188_/X _11330_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11331_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14050_ _14056_/CLK _14050_/D vssd1 vssd1 vccd1 vccd1 _14050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11262_ _11260_/Y _11213_/X _11261_/Y _11215_/X vssd1 vssd1 vccd1 vccd1 _11262_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13001_ _12580_/X _13000_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10213_ _11669_/A vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__buf_2
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11193_ _11429_/A vssd1 vssd1 vccd1 vccd1 _11193_/X sky130_fd_sc_hd__buf_2
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ _10146_/A _12424_/X vssd1 vssd1 vccd1 vccd1 _10144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10079_/A _10120_/A vssd1 vssd1 vccd1 vccd1 _12494_/S sky130_fd_sc_hd__or2_1
XFILLER_0_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _14139_/CLK _13903_/D vssd1 vssd1 vccd1 vccd1 _13903_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13834_ _14107_/CLK _13834_/D vssd1 vssd1 vccd1 vccd1 _13834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13765_ _14120_/CLK _13765_/D vssd1 vssd1 vccd1 vccd1 _13765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10977_ _11449_/A vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12716_ _09569_/X input332/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13696_ _14173_/CLK _13696_/D vssd1 vssd1 vccd1 vccd1 _13696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ _13337_/Q _12646_/X _12647_/S vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__mux2_1
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12578_ _13308_/Q _12577_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12578_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _14637_/CLK _14317_/D vssd1 vssd1 vccd1 vccd1 _14317_/Q sky130_fd_sc_hd__dfxtp_1
X_11529_ _13218_/Q _11485_/X _14041_/Q _11429_/X _11528_/X vssd1 vssd1 vccd1 vccd1
+ _11529_/X sky130_fd_sc_hd__a221o_4
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14248_ _14325_/CLK _14248_/D vssd1 vssd1 vccd1 vccd1 _14248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _14183_/CLK _14179_/D vssd1 vssd1 vccd1 vccd1 _14179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08740_ _13697_/Q _08677_/A _08579_/X _08679_/A _08737_/X vssd1 vssd1 vccd1 vccd1
+ _13697_/D sky130_fd_sc_hd__o221a_1
XFILLER_171_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08671_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08671_/X sky130_fd_sc_hd__buf_2
XFILLER_113_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _14250_/Q _07561_/A _07401_/X _07563_/A _07617_/X vssd1 vssd1 vccd1 vccd1
+ _14250_/D sky130_fd_sc_hd__o221a_1
XFILLER_199_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07553_ _14287_/Q _07488_/A _07480_/X _07490_/A _07550_/X vssd1 vssd1 vccd1 vccd1
+ _14287_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06504_ _06504_/A _06504_/B vssd1 vssd1 vccd1 vccd1 _06508_/A sky130_fd_sc_hd__or2_1
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _07484_/A _08340_/B _08744_/C _08091_/D vssd1 vssd1 vccd1 vccd1 _11679_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_74_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _13451_/Q _09215_/X _08914_/X _09217_/X _09219_/X vssd1 vssd1 vccd1 vccd1
+ _13451_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09154_ _13490_/Q _09146_/X _08914_/X _09148_/X _09149_/X vssd1 vssd1 vccd1 vccd1
+ _13490_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08105_ _08829_/A vssd1 vssd1 vccd1 vccd1 _08105_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09085_ _13529_/Q _09077_/X _08914_/X _09079_/X _09084_/X vssd1 vssd1 vccd1 vccd1
+ _13529_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08036_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 la_data_in[30] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_1
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__inv_2
XFILLER_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08938_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08938_/X sky130_fd_sc_hd__buf_2
XPHY_6214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _08869_/A vssd1 vssd1 vccd1 vccd1 _08869_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater680 _13368_/CLK vssd1 vssd1 vccd1 vccd1 _14071_/CLK sky130_fd_sc_hd__buf_12
X_10900_ _13553_/Q _10720_/X _13794_/Q _10721_/X vssd1 vssd1 vccd1 vccd1 _10900_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ _14127_/Q vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__inv_2
XPHY_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater691 _12619_/S vssd1 vssd1 vccd1 vccd1 _12647_/S sky130_fd_sc_hd__buf_6
XFILLER_166_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ _10826_/Y _10735_/X _10827_/Y _10737_/X _10830_/X vssd1 vssd1 vccd1 vccd1
+ _10838_/C sky130_fd_sc_hd__o221a_1
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _14120_/CLK _13550_/D vssd1 vssd1 vccd1 vccd1 _13550_/Q sky130_fd_sc_hd__dfxtp_1
X_10762_ _13394_/Q _10568_/X _13706_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _10762_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _12500_/X _06989_/X _12603_/S vssd1 vssd1 vccd1 vccd1 _12501_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _14595_/CLK _13481_/D vssd1 vssd1 vccd1 vccd1 _13481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10693_ _11403_/A vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12432_ _12431_/X _06897_/X _12603_/S vssd1 vssd1 vccd1 vccd1 _12432_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ _13201_/Q _12362_/X input78/X vssd1 vssd1 vccd1 vccd1 _12363_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14102_ _14110_/CLK _14102_/D vssd1 vssd1 vccd1 vccd1 _14102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11314_ _14076_/Q vssd1 vssd1 vccd1 vccd1 _11314_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12294_ _11590_/Y _14549_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12294_/X sky130_fd_sc_hd__mux2_4
XFILLER_120_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14033_ _14114_/CLK _14033_/D vssd1 vssd1 vccd1 vccd1 _14033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11245_ _13996_/Q vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11176_ _11412_/A vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10127_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _12443_/S sky130_fd_sc_hd__or2_1
XFILLER_114_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _12510_/X _10058_/B _10058_/C vssd1 vssd1 vccd1 vccd1 _10058_/Y sky130_fd_sc_hd__nor3_4
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13817_ _14130_/CLK _13817_/D vssd1 vssd1 vccd1 vccd1 _13817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13748_ _14121_/CLK _13748_/D vssd1 vssd1 vccd1 vccd1 _13748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _14146_/CLK _13679_/D vssd1 vssd1 vccd1 vccd1 _13679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09910_ _13312_/Q _09906_/Y _09912_/B vssd1 vssd1 vccd1 vccd1 _09910_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09841_ _09781_/A _09781_/B _09840_/Y vssd1 vssd1 vccd1 vccd1 _09841_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_193_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09772_ _09772_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__or2_1
X_06984_ _06991_/A _06984_/B vssd1 vssd1 vccd1 vccd1 _14566_/D sky130_fd_sc_hd__nor2_1
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08723_ _08723_/A vssd1 vssd1 vccd1 vccd1 _08723_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08654_ _13744_/Q _08588_/A _08577_/X _08591_/A _08653_/X vssd1 vssd1 vccd1 vccd1
+ _13744_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07605_ _07605_/A vssd1 vssd1 vccd1 vccd1 _07605_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08585_ _08745_/A _11648_/A vssd1 vssd1 vccd1 vccd1 _08644_/A sky130_fd_sc_hd__or2_2
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07536_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07536_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07467_ _07467_/A vssd1 vssd1 vccd1 vccd1 _07467_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09207_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07398_ _14369_/Q _07387_/X _07396_/X _07389_/X _07397_/X vssd1 vssd1 vccd1 vccd1
+ _14369_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09137_ _09137_/A vssd1 vssd1 vccd1 vccd1 _09137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09068_ _09120_/A vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__buf_2
XFILLER_178_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ _14053_/Q _07955_/A _07876_/X _07957_/A _08017_/X vssd1 vssd1 vccd1 vccd1
+ _14053_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _13477_/Q vssd1 vssd1 vccd1 vccd1 _11030_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12981_ _12570_/X _12980_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__mux2_1
XPHY_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11932_ _14401_/Q vssd1 vssd1 vccd1 vccd1 _11932_/Y sky130_fd_sc_hd__inv_2
XPHY_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _11861_/Y _11693_/X _11862_/Y _11695_/X vssd1 vssd1 vccd1 vccd1 _11863_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _14470_/CLK _13602_/D vssd1 vssd1 vccd1 vccd1 _13602_/Q sky130_fd_sc_hd__dfxtp_1
X_10814_ _13987_/Q vssd1 vssd1 vccd1 vccd1 _10814_/Y sky130_fd_sc_hd__inv_2
XPHY_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11792_/Y _11648_/X _11793_/Y _11650_/X vssd1 vssd1 vccd1 vccd1 _11794_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14582_ _14621_/CLK _14582_/D vssd1 vssd1 vccd1 vccd1 _14582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13533_ _14123_/CLK _13533_/D vssd1 vssd1 vccd1 vccd1 _13533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _11455_/A vssd1 vssd1 vccd1 vccd1 _10745_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13464_ _14173_/CLK _13464_/D vssd1 vssd1 vccd1 vccd1 _13464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _10674_/Y _10498_/X _10675_/Y _10501_/X vssd1 vssd1 vccd1 vccd1 _10676_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12415_ _12414_/X _13216_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13395_ _14183_/CLK _13395_/D vssd1 vssd1 vccd1 vccd1 _13395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12346_ _12345_/X _13191_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12346_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12277_ _12069_/Y _13378_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12277_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14016_ _14047_/CLK _14016_/D vssd1 vssd1 vccd1 vccd1 _14016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11228_ _11197_/X _11228_/B _11228_/C _11228_/D vssd1 vssd1 vccd1 vccd1 _11229_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_116_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11159_ _11159_/A _11159_/B _11159_/C _11159_/D vssd1 vssd1 vccd1 vccd1 _11159_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_81_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput280 la_oenb[87] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__buf_1
Xinput291 la_oenb[97] vssd1 vssd1 vccd1 vccd1 input291/X sky130_fd_sc_hd__buf_1
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _13882_/Q _08363_/X _08132_/X _08364_/X _08367_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/D sky130_fd_sc_hd__o221a_1
XFILLER_189_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07321_ _07387_/A vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07252_ _14436_/Q _07248_/X _06738_/X _07250_/X _07244_/X vssd1 vssd1 vccd1 vccd1
+ _14436_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07183_ _14473_/Q _07174_/X _06745_/X _07176_/X _07181_/X vssd1 vssd1 vccd1 vccd1
+ _14473_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09824_ _09824_/A vssd1 vssd1 vccd1 vccd1 _09824_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09755_ _13333_/Q vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__inv_2
X_06967_ _14570_/Q vssd1 vssd1 vccd1 vccd1 _06967_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08706_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08706_/X sky130_fd_sc_hd__clkbuf_2
X_09686_ _09682_/X _09685_/X _09682_/X _09685_/X vssd1 vssd1 vccd1 vccd1 _09686_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06898_ _06880_/X _12293_/X _06897_/X _06883_/X vssd1 vssd1 vccd1 vccd1 _06899_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08637_ _08637_/A vssd1 vssd1 vccd1 vccd1 _08637_/X sky130_fd_sc_hd__buf_1
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _13788_/Q _08565_/X _08566_/X _08567_/X _08563_/X vssd1 vssd1 vccd1 vccd1
+ _13788_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07519_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _08565_/A vssd1 vssd1 vccd1 vccd1 _08552_/A sky130_fd_sc_hd__buf_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10530_ _13864_/Q vssd1 vssd1 vccd1 vccd1 _10530_/Y sky130_fd_sc_hd__inv_2
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10461_ _11658_/A vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12200_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13180_ _14581_/Q _14582_/Q _14579_/Q _14580_/Q _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13180_/X sky130_fd_sc_hd__mux4_2
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10392_ _13862_/Q vssd1 vssd1 vccd1 vccd1 _10392_/Y sky130_fd_sc_hd__inv_2
X_12131_ vssd1 vssd1 vccd1 vccd1 _12131_/HI _12131_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _09791_/A _12057_/X _09903_/A _12058_/X vssd1 vssd1 vccd1 vccd1 _12062_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11013_ _11013_/A vssd1 vssd1 vccd1 vccd1 _11013_/X sky130_fd_sc_hd__buf_2
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12964_ _12562_/X input334/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12964_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _13419_/Q _11747_/X _13738_/Q _09601_/A _11914_/X vssd1 vssd1 vccd1 vccd1
+ _11948_/B sky130_fd_sc_hd__a221oi_2
XPHY_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12534_/X _12894_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__mux2_1
XPHY_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14634_ _14637_/CLK _14634_/D vssd1 vssd1 vccd1 vccd1 _14634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11846_ _13729_/Q _11642_/X _14048_/Q _11663_/X _11845_/X vssd1 vssd1 vccd1 vccd1
+ _11846_/X sky130_fd_sc_hd__a221o_2
XPHY_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11777_ _13493_/Q vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__inv_2
X_14565_ _14573_/CLK _14565_/D vssd1 vssd1 vccd1 vccd1 _14565_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10728_ _14609_/Q vssd1 vssd1 vccd1 vccd1 _10728_/Y sky130_fd_sc_hd__inv_2
X_13516_ _14110_/CLK _13516_/D vssd1 vssd1 vccd1 vccd1 _13516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14496_ _14621_/CLK _14496_/D vssd1 vssd1 vccd1 vccd1 _14496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10659_ _10657_/Y _10455_/X _10658_/Y _10458_/X vssd1 vssd1 vccd1 vccd1 _10659_/X
+ sky130_fd_sc_hd__o22a_1
X_13447_ _14183_/CLK _13447_/D vssd1 vssd1 vccd1 vccd1 _13447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13378_ _14538_/CLK _13378_/D vssd1 vssd1 vccd1 vccd1 _13378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12329_ _13196_/Q input94/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07870_ _14136_/Q _07863_/X _07790_/X _07864_/X _07865_/X vssd1 vssd1 vccd1 vccd1
+ _14136_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06821_ _07028_/A vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09540_ _09530_/X _09539_/X _13278_/Q _09531_/X vssd1 vssd1 vccd1 vccd1 _13246_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06752_ _08917_/A vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__buf_4
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09471_ _13282_/Q _09464_/X _12277_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _13282_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_168_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06683_ _06586_/A _06682_/Y _06586_/Y _06682_/A vssd1 vssd1 vccd1 vccd1 _06683_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08422_ _13854_/Q _08415_/X _08103_/X _08417_/X _08421_/X vssd1 vssd1 vccd1 vccd1
+ _13854_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08353_ _08396_/A vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07304_ _07558_/A _11675_/A vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__or2_2
X_08284_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08284_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07235_ _07558_/A _10165_/A vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__or2_2
XFILLER_34_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07166_ _07166_/A vssd1 vssd1 vccd1 vccd1 _07166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07097_ _14519_/Q _07092_/X _06714_/X _07094_/X _07096_/X vssd1 vssd1 vccd1 vccd1
+ _14519_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput540 _12168_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput551 _12178_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__clkbuf_2
Xoutput562 _12188_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput573 _12234_/X vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput584 _13272_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput595 _13282_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09807_ _13347_/Q vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__inv_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07999_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07999_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09738_ _10058_/C _12509_/S vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__or2_2
XFILLER_210_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09669_ _09667_/X _09668_/X _09667_/X _09668_/X vssd1 vssd1 vccd1 vccd1 _09669_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11700_ _14084_/Q vssd1 vssd1 vccd1 vccd1 _11700_/Y sky130_fd_sc_hd__inv_2
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _09589_/X input356/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__mux2_1
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B _11631_/C _11631_/D vssd1 vssd1 vccd1 vccd1 _11631_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _13847_/Q vssd1 vssd1 vccd1 vccd1 _11562_/Y sky130_fd_sc_hd__inv_2
X_14350_ _14629_/CLK _14350_/D vssd1 vssd1 vccd1 vccd1 _14350_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _14448_/Q vssd1 vssd1 vccd1 vccd1 _10513_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13301_ _13877_/CLK _13301_/D vssd1 vssd1 vccd1 vccd1 _13301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _14637_/CLK _14281_/D vssd1 vssd1 vccd1 vccd1 _14281_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _11488_/Y _11435_/X _11489_/Y _11437_/X _11492_/X vssd1 vssd1 vccd1 vccd1
+ _11506_/B sky130_fd_sc_hd__o221a_2
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13232_ _13352_/CLK _13232_/D vssd1 vssd1 vccd1 vccd1 _13264_/Q sky130_fd_sc_hd__dfxtp_2
X_10444_ _11646_/A vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _12659_/X _13162_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ _14134_/Q vssd1 vssd1 vccd1 vccd1 _10375_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ vssd1 vssd1 vccd1 vccd1 _12114_/HI _12114_/LO sky130_fd_sc_hd__conb_1
X_13094_ _13093_/X _12625_/X _13110_/S vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12045_ _09778_/A _12043_/X _09890_/A _12044_/X vssd1 vssd1 vccd1 vccd1 _12045_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_26_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13996_ _13996_/CLK _13996_/D vssd1 vssd1 vccd1 vccd1 _13996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12947_ _12553_/X _12946_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_160 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12530_/X _12877_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _06603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_182 input335/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_193 input356/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14617_ _14627_/CLK _14617_/D vssd1 vssd1 vccd1 vccd1 _14617_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _11824_/Y _11633_/X _11825_/Y _11635_/X _11828_/X vssd1 vssd1 vccd1 vccd1
+ _11866_/A sky130_fd_sc_hd__o221a_2
XFILLER_18_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _14611_/CLK _14548_/D vssd1 vssd1 vccd1 vccd1 _14548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14479_ _14481_/CLK _14479_/D vssd1 vssd1 vccd1 vccd1 _14479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07020_ _14558_/Q _07014_/X _06714_/X _07017_/X _07018_/X vssd1 vssd1 vccd1 vccd1
+ _14558_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08971_ _08971_/A vssd1 vssd1 vccd1 vccd1 _08971_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07922_ _14109_/Q _07918_/X _07762_/X _07919_/X _07921_/X vssd1 vssd1 vccd1 vccd1
+ _14109_/D sky130_fd_sc_hd__o221a_1
XFILLER_155_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07853_ _14146_/Q _07845_/X _07852_/X _07846_/X _07848_/X vssd1 vssd1 vccd1 vccd1
+ _14146_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06804_ _14613_/Q _06787_/X _06801_/X _06790_/X _06803_/X vssd1 vssd1 vccd1 vccd1
+ _14613_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _08175_/A vssd1 vssd1 vccd1 vccd1 _07784_/X sky130_fd_sc_hd__buf_4
XFILLER_186_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06735_ _07719_/A vssd1 vssd1 vccd1 vccd1 _06735_/X sky130_fd_sc_hd__buf_2
X_09523_ _09514_/X _09522_/X _13284_/Q _09517_/X vssd1 vssd1 vccd1 vccd1 _13252_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ _09456_/A _12943_/X vssd1 vssd1 vccd1 vccd1 _13290_/D sky130_fd_sc_hd__and2_1
X_06666_ _06634_/X _06665_/X _06634_/X _06665_/X vssd1 vssd1 vccd1 vccd1 _06666_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ _13860_/Q _08344_/A _08188_/X _08346_/A _08400_/X vssd1 vssd1 vccd1 vccd1
+ _13860_/D sky130_fd_sc_hd__o221a_1
X_09385_ _09388_/A _13167_/X vssd1 vssd1 vccd1 vccd1 _13346_/D sky130_fd_sc_hd__and2_1
XFILLER_90_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06597_ _06593_/Y _08935_/A _08914_/A _06596_/Y vssd1 vssd1 vccd1 vccd1 _06598_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08336_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08336_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08267_ _13937_/Q _08198_/A _08190_/X _08201_/A _08264_/X vssd1 vssd1 vccd1 vccd1
+ _13937_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _07218_/A vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08198_ _08198_/A vssd1 vssd1 vccd1 vccd1 _08198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07149_ _14488_/Q _07144_/X _06831_/X _07145_/X _07147_/X vssd1 vssd1 vccd1 vccd1
+ _14488_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10160_ _10154_/Y _10156_/X _10157_/Y _10159_/X vssd1 vssd1 vccd1 vccd1 _10160_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput370 _12207_/X vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput381 _12217_/X vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput392 _12227_/X vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10091_ _10094_/A _12484_/X vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__nor2_8
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13850_ _14094_/CLK _13850_/D vssd1 vssd1 vccd1 vccd1 _13850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _12512_/X _12800_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12801_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ _14123_/CLK _13781_/D vssd1 vssd1 vccd1 vccd1 _13781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10993_ _10993_/A _10993_/B _10993_/C _10993_/D vssd1 vssd1 vccd1 vccd1 _10993_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_210_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12732_ _09539_/X input345/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12732_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _13345_/Q _12662_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__mux2_1
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14402_ _14633_/CLK _14402_/D vssd1 vssd1 vccd1 vccd1 _14402_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11614_ _14628_/Q vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__inv_2
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12594_ _13316_/Q _12593_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12594_/X sky130_fd_sc_hd__mux2_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14333_ _14527_/CLK _14333_/D vssd1 vssd1 vccd1 vccd1 _14333_/Q sky130_fd_sc_hd__dfxtp_1
X_11545_ _14470_/Q vssd1 vssd1 vccd1 vccd1 _11545_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11476_ _13884_/Q vssd1 vssd1 vccd1 vccd1 _11476_/Y sky130_fd_sc_hd__inv_2
X_14264_ _14305_/CLK _14264_/D vssd1 vssd1 vccd1 vccd1 _14264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10427_ _11635_/A vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__buf_4
X_13215_ _14459_/CLK _13215_/D vssd1 vssd1 vccd1 vccd1 _13215_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_193_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14195_ _14529_/CLK _14195_/D vssd1 vssd1 vccd1 vccd1 _14195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10358_ _10356_/Y _10195_/X _10357_/Y _10198_/X vssd1 vssd1 vccd1 vccd1 _10358_/X
+ sky130_fd_sc_hd__o22a_1
X_13146_ _13145_/X _12651_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13077_ _12618_/X _13076_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10289_ _10287_/Y _10234_/X _10288_/Y _10237_/X vssd1 vssd1 vccd1 vccd1 _10289_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12028_ _12023_/Y _10242_/A _12024_/Y _10245_/A _12027_/X vssd1 vssd1 vccd1 vccd1
+ _12029_/D sky130_fd_sc_hd__o221a_1
XFILLER_152_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13979_ _14100_/CLK _13979_/D vssd1 vssd1 vccd1 vccd1 _13979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06520_ _09272_/A vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09170_ _13480_/Q _09163_/X _08942_/X _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1
+ _13480_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08121_ _14004_/Q _08109_/X _08119_/X _08112_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _14004_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _14038_/Q _08045_/X _07742_/X _08046_/X _08050_/X vssd1 vssd1 vccd1 vccd1
+ _14038_/D sky130_fd_sc_hd__o221a_1
X_07003_ _06857_/A _12322_/X _10057_/A _06861_/A vssd1 vssd1 vccd1 vccd1 _07004_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput109 la_data_in[48] vssd1 vssd1 vccd1 vccd1 _06596_/A sky130_fd_sc_hd__clkbuf_2
X_08954_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08954_/X sky130_fd_sc_hd__buf_4
XFILLER_9_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07905_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08885_ _13620_/Q _08818_/A _08577_/X _08820_/A _08880_/X vssd1 vssd1 vccd1 vccd1
+ _13620_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ _14155_/Q _07829_/X _07742_/X _07830_/X _07831_/X vssd1 vssd1 vccd1 vccd1
+ _14155_/D sky130_fd_sc_hd__o221a_1
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07767_ _08158_/A vssd1 vssd1 vccd1 vccd1 _07767_/X sky130_fd_sc_hd__buf_4
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09506_ _13257_/Q _09500_/X _12252_/X _09501_/X vssd1 vssd1 vccd1 vccd1 _13257_/D
+ sky130_fd_sc_hd__o22a_1
X_06718_ _08825_/A vssd1 vssd1 vccd1 vccd1 _07710_/A sky130_fd_sc_hd__clkbuf_4
X_07698_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09438_/A _13015_/X vssd1 vssd1 vccd1 vccd1 _13304_/D sky130_fd_sc_hd__and2_1
X_06649_ _06644_/X _06648_/X _06644_/X _06648_/X vssd1 vssd1 vccd1 vccd1 _06649_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09368_ _09370_/A _12855_/X vssd1 vssd1 vccd1 vccd1 _13360_/D sky130_fd_sc_hd__and2_1
XFILLER_178_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08319_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ _13409_/Q _09294_/X _08128_/A _09295_/X _09298_/X vssd1 vssd1 vccd1 vccd1
+ _13409_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_60 _07788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_71 _08165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _08336_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11330_ _13523_/Q vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_93 _08935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ _14269_/Q vssd1 vssd1 vccd1 vccd1 _11261_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _14482_/Q vssd1 vssd1 vccd1 vccd1 _10212_/Y sky130_fd_sc_hd__inv_2
X_13000_ _12580_/X input342/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13000_/X sky130_fd_sc_hd__mux2_1
X_11192_ _11175_/Y _11176_/X _11181_/X _11186_/X _11191_/X vssd1 vssd1 vccd1 vccd1
+ _11229_/C sky130_fd_sc_hd__o2111a_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _10143_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _12422_/S sky130_fd_sc_hd__or2_1
XFILLER_66_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10074_ _10098_/A _10113_/A vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__or2_1
XPHY_6930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _14139_/CLK _13902_/D vssd1 vssd1 vccd1 vccd1 _13902_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13833_ _14107_/CLK _13833_/D vssd1 vssd1 vccd1 vccd1 _13833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13764_ _13996_/CLK _13764_/D vssd1 vssd1 vccd1 vccd1 _13764_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _14185_/Q vssd1 vssd1 vccd1 vccd1 _10976_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12715_ _09567_/X _12714_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13203_/D sky130_fd_sc_hd__mux2_1
X_13695_ _14173_/CLK _13695_/D vssd1 vssd1 vccd1 vccd1 _13695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12646_ _09825_/Y _13337_/Q _12650_/S vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__mux2_1
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ _09939_/X _13308_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__mux2_1
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14316_ _14527_/CLK _14316_/D vssd1 vssd1 vccd1 vccd1 _14316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _13566_/Q _11430_/X _13807_/Q _11431_/X vssd1 vssd1 vccd1 vccd1 _11528_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14247_ _14325_/CLK _14247_/D vssd1 vssd1 vccd1 vccd1 _14247_/Q sky130_fd_sc_hd__dfxtp_1
X_11459_ _11459_/A vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14178_ _14178_/CLK _14178_/D vssd1 vssd1 vccd1 vccd1 _14178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13129_ _12643_/X _13128_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08670_ _13735_/Q _08662_/A _08501_/X _08663_/A _08665_/X vssd1 vssd1 vccd1 vccd1
+ _13735_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07621_ _14251_/Q _07561_/A _07399_/X _07563_/A _07617_/X vssd1 vssd1 vccd1 vccd1
+ _14251_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07552_ _14288_/Q _07488_/A _07403_/X _07490_/A _07550_/X vssd1 vssd1 vccd1 vccd1
+ _14288_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06503_ _06503_/A _06503_/B _06503_/C _06503_/D vssd1 vssd1 vccd1 vccd1 _06504_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_59_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07483_ _08482_/D vssd1 vssd1 vccd1 vccd1 _08091_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _13452_/Q _09215_/X _08912_/X _09217_/X _09219_/X vssd1 vssd1 vccd1 vccd1
+ _13452_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09153_ _13491_/Q _09146_/X _08912_/X _09148_/X _09149_/X vssd1 vssd1 vccd1 vccd1
+ _13491_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08104_ _14010_/Q _08095_/X _08103_/X _08097_/X _08089_/X vssd1 vssd1 vccd1 vccd1
+ _14010_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09084_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08035_ _08078_/A vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__buf_2
Xinput80 la_data_in[21] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_1
XFILLER_200_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput91 la_data_in[31] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_1
XFILLER_66_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09986_ _13364_/Q _09986_/B vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ _09138_/A vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__buf_2
XPHY_6215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _08868_/A vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater670 _14143_/CLK vssd1 vssd1 vccd1 vccd1 _14183_/CLK sky130_fd_sc_hd__buf_12
XFILLER_6_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07819_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater681 _13368_/CLK vssd1 vssd1 vccd1 vccd1 _13352_/CLK sky130_fd_sc_hd__buf_12
XPHY_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater692 _12651_/S vssd1 vssd1 vccd1 vccd1 _12619_/S sky130_fd_sc_hd__buf_8
XPHY_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08799_ _13665_/Q _08792_/X _08562_/X _08793_/X _08794_/X vssd1 vssd1 vccd1 vccd1
+ _13665_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10830_ _10828_/Y _10739_/X _10829_/Y _10741_/X vssd1 vssd1 vccd1 vccd1 _10830_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10761_ _10756_/Y _10687_/X _10757_/Y _10689_/X _10760_/X vssd1 vssd1 vccd1 vccd1
+ _10797_/A sky130_fd_sc_hd__o221a_2
XFILLER_0_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _12509_/X _06989_/X _12500_/S vssd1 vssd1 vccd1 vccd1 _12500_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10692_ _13627_/Q vssd1 vssd1 vccd1 vccd1 _10692_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13480_ _14595_/CLK _13480_/D vssd1 vssd1 vccd1 vccd1 _13480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12509_/X _06897_/X _12431_/S vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12362_ _13201_/Q input98/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14101_ _14110_/CLK _14101_/D vssd1 vssd1 vccd1 vccd1 _14101_/Q sky130_fd_sc_hd__dfxtp_1
X_11313_ _11313_/A _11313_/B _11313_/C _11313_/D vssd1 vssd1 vccd1 vccd1 _11313_/Y
+ sky130_fd_sc_hd__nand4_4
X_12293_ _11631_/Y _14550_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__mux2_2
XFILLER_120_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14032_ _14119_/CLK _14032_/D vssd1 vssd1 vccd1 vccd1 _14032_/Q sky130_fd_sc_hd__dfxtp_1
X_11244_ _11242_/Y _11183_/X _11243_/Y _11185_/X vssd1 vssd1 vccd1 vccd1 _11244_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11175_ _13956_/Q vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10126_ _10126_/A _12448_/X vssd1 vssd1 vccd1 vccd1 _10126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10057_ _10057_/A _10060_/A vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13816_ _14130_/CLK _13816_/D vssd1 vssd1 vccd1 vccd1 _13816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13747_ _14094_/CLK _13747_/D vssd1 vssd1 vccd1 vccd1 _13747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10959_ _11431_/A vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13678_ _14146_/CLK _13678_/D vssd1 vssd1 vccd1 vccd1 _13678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12629_ _13330_/Q _12628_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__mux2_1
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _09840_/A vssd1 vssd1 vccd1 vccd1 _09840_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09771_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__or2_1
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06983_ _06974_/X _12316_/X _06982_/Y _06976_/X vssd1 vssd1 vccd1 vccd1 _06984_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08722_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08653_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08653_/X sky130_fd_sc_hd__clkbuf_4
XPHY_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07604_ _14262_/Q _07597_/X _07370_/X _07598_/X _07601_/X vssd1 vssd1 vccd1 vccd1
+ _14262_/D sky130_fd_sc_hd__o221a_1
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08584_ _08744_/A _09201_/B _08584_/C _08584_/D vssd1 vssd1 vccd1 vccd1 _11648_/A
+ sky130_fd_sc_hd__or4_4
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07535_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07466_ _14335_/Q _07459_/X _07383_/X _07460_/X _07461_/X vssd1 vssd1 vccd1 vccd1
+ _14335_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09205_ _09205_/A vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__clkbuf_2
X_07397_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07397_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09136_ _09189_/A vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09067_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ _14054_/Q _07955_/A _07800_/X _07957_/A _08017_/X vssd1 vssd1 vccd1 vccd1
+ _14054_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09969_ _09969_/A vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__inv_2
XPHY_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _12570_/X input361/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11931_ _14635_/Q vssd1 vssd1 vccd1 vccd1 _11931_/Y sky130_fd_sc_hd__inv_2
XPHY_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _14477_/Q vssd1 vssd1 vccd1 vccd1 _11862_/Y sky130_fd_sc_hd__inv_2
XPHY_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13601_ _14305_/CLK _13601_/D vssd1 vssd1 vccd1 vccd1 _13601_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _10811_/Y _10709_/X _10812_/Y _10711_/X vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_183_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14581_ _14621_/CLK _14581_/D vssd1 vssd1 vccd1 vccd1 _14581_/Q sky130_fd_sc_hd__dfxtp_2
X_11793_ _13891_/Q vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__inv_2
XPHY_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13532_ _14123_/CLK _13532_/D vssd1 vssd1 vccd1 vccd1 _13532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10744_ _13907_/Q vssd1 vssd1 vccd1 vccd1 _10744_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13463_ _14173_/CLK _13463_/D vssd1 vssd1 vccd1 vccd1 _13463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10675_ _14257_/Q vssd1 vssd1 vccd1 vccd1 _10675_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12414_ _13216_/Q _12413_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12414_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13394_ _14183_/CLK _13394_/D vssd1 vssd1 vccd1 vccd1 _13394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12345_ _13191_/Q _12344_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12345_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12276_ _12068_/Y _13377_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14015_ _14047_/CLK _14015_/D vssd1 vssd1 vccd1 vccd1 _14015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11227_ _11218_/Y _11219_/X _11220_/Y _11221_/X _11226_/X vssd1 vssd1 vccd1 vccd1
+ _11228_/D sky130_fd_sc_hd__o221a_1
XFILLER_68_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11158_ _11139_/X _11158_/B _11158_/C _11158_/D vssd1 vssd1 vccd1 vccd1 _11159_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ _10114_/A _12469_/X vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11089_ _11087_/Y _10942_/X _11088_/Y _10944_/X vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput270 la_oenb[78] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__buf_1
XFILLER_42_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput281 la_oenb[88] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_hd__buf_1
XFILLER_42_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput292 la_oenb[98] vssd1 vssd1 vccd1 vccd1 input292/X sky130_fd_sc_hd__buf_1
XFILLER_23_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07320_ _14399_/Q _07307_/X _07317_/X _07309_/X _07319_/X vssd1 vssd1 vccd1 vccd1
+ _14399_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07251_ _14437_/Q _07248_/X _06735_/X _07250_/X _07244_/X vssd1 vssd1 vccd1 vccd1
+ _14437_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07182_ _14474_/Q _07174_/X _07031_/X _07176_/X _07181_/X vssd1 vssd1 vccd1 vccd1
+ _14474_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _13336_/Q _09820_/Y _09787_/B vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _13334_/Q vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__inv_2
X_06966_ _06972_/A _06966_/B vssd1 vssd1 vccd1 vccd1 _14571_/D sky130_fd_sc_hd__nor2_1
XFILLER_210_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08705_ _13719_/Q _08698_/X _08523_/X _08699_/X _08704_/X vssd1 vssd1 vccd1 vccd1
+ _13719_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09685_ _09668_/X _09684_/Y _09668_/X _09684_/Y vssd1 vssd1 vccd1 vccd1 _09685_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06897_ _06897_/A vssd1 vssd1 vccd1 vccd1 _06897_/X sky130_fd_sc_hd__clkbuf_4
X_08636_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08636_/X sky130_fd_sc_hd__buf_1
XFILLER_110_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08567_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07518_ _14310_/Q _07516_/X _07349_/X _07517_/X _07511_/X vssd1 vssd1 vccd1 vccd1
+ _14310_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08498_ _13814_/Q _08486_/X _08496_/X _08488_/X _08497_/X vssd1 vssd1 vccd1 vccd1
+ _13814_/D sky130_fd_sc_hd__o221a_1
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _14345_/Q _07440_/X _07358_/X _07441_/X _07444_/X vssd1 vssd1 vccd1 vccd1
+ _14345_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10460_ _13980_/Q vssd1 vssd1 vccd1 vccd1 _10460_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _09119_/A vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__clkbuf_2
X_10391_ _13745_/Q vssd1 vssd1 vccd1 vccd1 _10391_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ vssd1 vssd1 vccd1 vccd1 _12130_/HI _12130_/LO sky130_fd_sc_hd__conb_1
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12061_ _09790_/A _12057_/X _09902_/A _12058_/X vssd1 vssd1 vccd1 vccd1 _12061_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_78_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _11002_/Y _10940_/X _11005_/X _11008_/X _11011_/X vssd1 vssd1 vccd1 vccd1
+ _11035_/C sky130_fd_sc_hd__o2111a_4
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _12560_/X _12962_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12963_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11914_ _14245_/Q _11830_/X _14440_/Q _11831_/X vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _12534_/X _12893_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12894_/X sky130_fd_sc_hd__mux2_1
XPHY_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/CLK _14633_/D vssd1 vssd1 vccd1 vccd1 _14633_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _13573_/Q _11664_/X _13814_/Q _11665_/X vssd1 vssd1 vccd1 vccd1 _11845_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14573_/CLK _14564_/D vssd1 vssd1 vccd1 vccd1 _14564_/Q sky130_fd_sc_hd__dfxtp_2
X_11776_ _14163_/Q vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13996_/CLK _13515_/D vssd1 vssd1 vccd1 vccd1 _13515_/Q sky130_fd_sc_hd__dfxtp_1
X_10727_ _11437_/A vssd1 vssd1 vccd1 vccd1 _10727_/X sky130_fd_sc_hd__buf_2
X_14495_ _14495_/CLK _14495_/D vssd1 vssd1 vccd1 vccd1 _14495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13446_ _14183_/CLK _13446_/D vssd1 vssd1 vccd1 vccd1 _13446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10658_ _14101_/Q vssd1 vssd1 vccd1 vccd1 _10658_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13377_ _14573_/CLK _13377_/D vssd1 vssd1 vccd1 vccd1 _13377_/Q sky130_fd_sc_hd__dfxtp_1
X_10589_ _10584_/Y _10478_/X _10585_/Y _10481_/X _10588_/X vssd1 vssd1 vccd1 vccd1
+ _10602_/B sky130_fd_sc_hd__o221a_2
XFILLER_182_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12328_ _12327_/X _13197_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12328_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12259_ _12045_/Y _13360_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06820_ _08171_/A vssd1 vssd1 vccd1 vccd1 _06820_/X sky130_fd_sc_hd__buf_2
XFILLER_116_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09470_ _13283_/Q _09464_/X _12278_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _13283_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06682_ _06682_/A vssd1 vssd1 vccd1 vccd1 _06682_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08421_ _08421_/A vssd1 vssd1 vccd1 vccd1 _08421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08352_ _13892_/Q _08344_/X _08105_/X _08346_/X _08349_/X vssd1 vssd1 vccd1 vccd1
+ _13892_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07303_ _08744_/A _09271_/B _09131_/C _09271_/D vssd1 vssd1 vccd1 vccd1 _11675_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_127_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08283_ _08326_/A vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_127_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07234_ _07484_/A _07878_/B _08744_/C _07630_/D vssd1 vssd1 vccd1 vccd1 _10165_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07165_ _07218_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07096_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07096_/X sky130_fd_sc_hd__buf_2
XFILLER_69_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput530 _12104_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput541 _12105_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput552 _12106_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput563 _12107_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput574 _12108_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput585 _13273_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput596 _13283_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09806_ _13346_/Q _09802_/Y _09808_/B vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07998_ _14067_/Q _07991_/X _07767_/X _07992_/X _07995_/X vssd1 vssd1 vccd1 vccd1
+ _14067_/D sky130_fd_sc_hd__o221a_1
XFILLER_169_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09737_ _12508_/S vssd1 vssd1 vccd1 vccd1 _10058_/C sky130_fd_sc_hd__inv_2
XFILLER_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06949_ _14575_/Q vssd1 vssd1 vccd1 vccd1 _06949_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ _14566_/Q _14565_/Q _06982_/Y _06985_/Y vssd1 vssd1 vccd1 vccd1 _09668_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08619_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08619_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09599_ _09599_/A vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__inv_2
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11630_ _11611_/X _11630_/B _11630_/C _11630_/D vssd1 vssd1 vccd1 vccd1 _11631_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11561_ _11559_/Y _11414_/X _11560_/Y _11416_/X vssd1 vssd1 vccd1 vccd1 _11561_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _13877_/CLK _13300_/D vssd1 vssd1 vccd1 vccd1 _13300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10512_ _11459_/A vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _14637_/CLK _14280_/D vssd1 vssd1 vccd1 vccd1 _14280_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11492_ _11490_/Y _11439_/X _11491_/Y _11441_/X vssd1 vssd1 vccd1 vccd1 _11492_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _13352_/CLK _13231_/D vssd1 vssd1 vccd1 vccd1 _13263_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10443_ _13941_/Q vssd1 vssd1 vccd1 vccd1 _10443_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13162_ _13161_/X _12659_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10374_ _13900_/Q vssd1 vssd1 vccd1 vccd1 _10374_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12113_ vssd1 vssd1 vccd1 vccd1 _12113_/HI _12113_/LO sky130_fd_sc_hd__conb_1
X_13093_ _12625_/X _13092_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12044_ _12065_/A vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__buf_2
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13995_ _13996_/CLK _13995_/D vssd1 vssd1 vccd1 vccd1 _13995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12946_ _12945_/X _12553_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_150 _11611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _12530_/X _12876_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__mux2_1
XANTENNA_161 _11969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 input330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14616_ _14627_/CLK _14616_/D vssd1 vssd1 vccd1 vccd1 _14616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ _11826_/Y _11637_/X _11827_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _11828_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_183 input336/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_194 input357/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14547_ _14611_/CLK _14547_/D vssd1 vssd1 vccd1 vccd1 _14547_/Q sky130_fd_sc_hd__dfxtp_1
X_11759_ _11757_/Y _11658_/X _11758_/Y _11660_/X vssd1 vssd1 vccd1 vccd1 _11759_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14478_ _14481_/CLK _14478_/D vssd1 vssd1 vccd1 vccd1 _14478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13429_ _14139_/CLK _13429_/D vssd1 vssd1 vccd1 vccd1 _13429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08970_ input96/X vssd1 vssd1 vccd1 vccd1 _08970_/X sky130_fd_sc_hd__buf_4
XFILLER_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07921_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07852_ _08243_/A vssd1 vssd1 vccd1 vccd1 _07852_/X sky130_fd_sc_hd__buf_4
XFILLER_211_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06803_ _07028_/A vssd1 vssd1 vccd1 vccd1 _06803_/X sky130_fd_sc_hd__clkbuf_2
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_110_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07783_ _07783_/A vssd1 vssd1 vccd1 vccd1 _07783_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _09533_/A _12403_/X vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__and2_1
XFILLER_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06734_ _08833_/A vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__buf_2
XFILLER_209_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09453_ _09456_/A _12939_/X vssd1 vssd1 vccd1 vccd1 _13291_/D sky130_fd_sc_hd__and2_1
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06665_ _08920_/A _08942_/A _06625_/Y _06614_/Y vssd1 vssd1 vccd1 vccd1 _06665_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _13861_/Q _08344_/A _08186_/X _08346_/A _08400_/X vssd1 vssd1 vccd1 vccd1
+ _13861_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09384_ _09388_/A _13163_/X vssd1 vssd1 vccd1 vccd1 _13347_/D sky130_fd_sc_hd__and2_1
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06596_ _06596_/A vssd1 vssd1 vccd1 vccd1 _06596_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08335_ _08383_/A vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08266_ _13938_/Q _08198_/A _08188_/X _08201_/A _08264_/X vssd1 vssd1 vccd1 vccd1
+ _13938_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07217_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07217_/X sky130_fd_sc_hd__clkbuf_2
X_08197_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07148_ _14489_/Q _07144_/X _07073_/X _07145_/X _07147_/X vssd1 vssd1 vccd1 vccd1
+ _14489_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput371 _12208_/X vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput382 _12218_/X vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10090_ _10090_/A _10132_/A vssd1 vssd1 vccd1 vccd1 _12482_/S sky130_fd_sc_hd__or2_1
XFILLER_82_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput393 _12228_/X vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ _12512_/X input358/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _14123_/CLK _13780_/D vssd1 vssd1 vccd1 vccd1 _13780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10992_ _10961_/X _10992_/B _10992_/C _10992_/D vssd1 vssd1 vccd1 vccd1 _10993_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_186_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12731_ _09578_/X _12730_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13199_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _09803_/Y _13345_/Q _12666_/S vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__mux2_1
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14401_ _14633_/CLK _14401_/D vssd1 vssd1 vccd1 vccd1 _14401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11613_ _14355_/Q vssd1 vssd1 vccd1 vccd1 _11613_/Y sky130_fd_sc_hd__inv_2
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _09924_/X _13316_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12593_/X sky130_fd_sc_hd__mux2_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _14527_/CLK _14332_/D vssd1 vssd1 vccd1 vccd1 _14332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _13488_/Q vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _14305_/CLK _14263_/D vssd1 vssd1 vccd1 vccd1 _14263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _13767_/Q vssd1 vssd1 vccd1 vccd1 _11475_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13214_ _14459_/CLK _13214_/D vssd1 vssd1 vccd1 vccd1 _13214_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ _13427_/Q vssd1 vssd1 vccd1 vccd1 _10426_/Y sky130_fd_sc_hd__inv_2
X_14194_ _14470_/CLK _14194_/D vssd1 vssd1 vccd1 vccd1 _14194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _12651_/X _13144_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10357_ _13503_/Q vssd1 vssd1 vccd1 vccd1 _10357_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13076_ _12618_/X input341/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10288_ _14249_/Q vssd1 vssd1 vccd1 vccd1 _10288_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12027_ _12025_/Y _10248_/A _12026_/Y _10251_/A vssd1 vssd1 vccd1 vccd1 _12027_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13978_ _14095_/CLK _13978_/D vssd1 vssd1 vccd1 vccd1 _13978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12929_ _12545_/X _12928_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08120_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08051_ _14039_/Q _08045_/X _07740_/X _08046_/X _08050_/X vssd1 vssd1 vccd1 vccd1
+ _14039_/D sky130_fd_sc_hd__o221a_1
XFILLER_102_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07002_ _14560_/Q vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__inv_2
XFILLER_50_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08953_ _13593_/Q _08944_/X _08632_/X _08946_/X _08951_/X vssd1 vssd1 vccd1 vccd1
+ _13593_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07904_ _14120_/Q _07902_/X _07733_/X _07903_/X _07897_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08884_ _13621_/Q _08876_/X _08574_/X _08877_/X _08880_/X vssd1 vssd1 vccd1 vccd1
+ _13621_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07835_ _14156_/Q _07829_/X _07740_/X _07830_/X _07831_/X vssd1 vssd1 vccd1 vccd1
+ _14156_/D sky130_fd_sc_hd__o221a_1
XFILLER_79_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07766_ _14185_/Q _07758_/X _07456_/X _07760_/X _07756_/X vssd1 vssd1 vccd1 vccd1
+ _14185_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _13258_/Q _09500_/X _12253_/X _09501_/X vssd1 vssd1 vccd1 vccd1 _13258_/D
+ sky130_fd_sc_hd__o22a_1
X_06717_ _14636_/Q _06530_/X _06714_/X _06716_/X _06723_/C1 vssd1 vssd1 vccd1 vccd1
+ _14636_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _14210_/Q _07634_/A _07403_/X _07636_/A _07692_/X vssd1 vssd1 vccd1 vccd1
+ _14210_/D sky130_fd_sc_hd__o221a_1
XFILLER_77_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09436_ _09438_/A _13011_/X vssd1 vssd1 vccd1 vccd1 _13305_/D sky130_fd_sc_hd__and2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06648_ _06646_/X _06647_/X _06646_/X _06647_/X vssd1 vssd1 vccd1 vccd1 _06648_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09367_ _09370_/A _12851_/X vssd1 vssd1 vccd1 vccd1 _13361_/D sky130_fd_sc_hd__and2_1
XFILLER_107_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06579_ _06573_/X _06578_/X _06573_/X _06578_/X vssd1 vssd1 vccd1 vccd1 _06579_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08318_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08318_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_50 _07719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09298_/X sky130_fd_sc_hd__buf_2
XANTENNA_61 _07792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_72 _08165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 _08480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _08288_/A vssd1 vssd1 vccd1 vccd1 _08249_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_94 _08940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11260_ _14191_/Q vssd1 vssd1 vccd1 vccd1 _11260_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _13191_/Q _09601_/A _14014_/Q _10203_/X _10210_/X vssd1 vssd1 vccd1 vccd1
+ _10211_/X sky130_fd_sc_hd__a221o_2
XFILLER_101_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ _11187_/Y _11188_/X _11189_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11191_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_161_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10146_/A _12427_/X vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10073_ _10080_/A _12499_/X vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__nor2_8
XFILLER_47_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _14139_/CLK _13901_/D vssd1 vssd1 vccd1 vccd1 _13901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13832_ _14107_/CLK _13832_/D vssd1 vssd1 vccd1 vccd1 _13832_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13763_ _13996_/CLK _13763_/D vssd1 vssd1 vccd1 vccd1 _13763_/Q sky130_fd_sc_hd__dfxtp_1
X_10975_ _11447_/A vssd1 vssd1 vccd1 vccd1 _10975_/X sky130_fd_sc_hd__buf_1
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _09567_/X _12713_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13694_ _14056_/CLK _13694_/D vssd1 vssd1 vccd1 vccd1 _13694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12645_ _13338_/Q _12644_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__mux2_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12576_ _13309_/Q _12575_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__mux2_1
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _14527_/CLK _14315_/D vssd1 vssd1 vccd1 vccd1 _14315_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11517_/Y _11412_/X _11520_/X _11523_/X _11526_/X vssd1 vssd1 vccd1 vccd1
+ _11549_/C sky130_fd_sc_hd__o2111a_4
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14246_ _14325_/CLK _14246_/D vssd1 vssd1 vccd1 vccd1 _14246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ _13486_/Q vssd1 vssd1 vccd1 vccd1 _11458_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10409_ _14291_/Q vssd1 vssd1 vccd1 vccd1 _10409_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14177_ _14529_/CLK _14177_/D vssd1 vssd1 vccd1 vccd1 _14177_/Q sky130_fd_sc_hd__dfxtp_1
X_11389_ _14155_/Q vssd1 vssd1 vccd1 vccd1 _11389_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13128_ _12643_/X input342/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13128_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13059_ _12608_/X _13058_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07620_ _14252_/Q _07613_/X _07396_/X _07614_/X _07617_/X vssd1 vssd1 vccd1 vccd1
+ _14252_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ _14289_/Q _07488_/A _07401_/X _07490_/A _07550_/X vssd1 vssd1 vccd1 vccd1
+ _14289_/D sky130_fd_sc_hd__o221a_1
XFILLER_4_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06502_ _06502_/A _06502_/B _06502_/C _06502_/D vssd1 vssd1 vccd1 vccd1 _06504_/A
+ sky130_fd_sc_hd__or4_4
X_07482_ _08989_/D vssd1 vssd1 vccd1 vccd1 _08482_/D sky130_fd_sc_hd__inv_2
XFILLER_62_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09221_ _13453_/Q _09215_/X _09009_/X _09217_/X _09219_/X vssd1 vssd1 vccd1 vccd1
+ _13453_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09152_ _13492_/Q _09146_/X _09009_/X _09148_/X _09149_/X vssd1 vssd1 vccd1 vccd1
+ _13492_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08103_ _08827_/A vssd1 vssd1 vccd1 vccd1 _08103_/X sky130_fd_sc_hd__buf_4
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09083_ _13530_/Q _09077_/X _08912_/X _09079_/X _09074_/X vssd1 vssd1 vccd1 vccd1
+ _13530_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08034_ _14048_/Q _08025_/X _07714_/X _08027_/X _08032_/X vssd1 vssd1 vccd1 vccd1
+ _14048_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput70 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
XFILLER_200_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput81 la_data_in[22] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_1
Xinput92 la_data_in[32] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _09985_/A vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__inv_2
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08936_ _08936_/A vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08867_ _13631_/Q _08860_/X _08549_/X _08861_/X _08863_/X vssd1 vssd1 vccd1 vccd1
+ _13631_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater660 _14047_/CLK vssd1 vssd1 vccd1 vccd1 _14056_/CLK sky130_fd_sc_hd__buf_8
XPHY_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ _07863_/A vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__buf_6
Xrepeater671 _14143_/CLK vssd1 vssd1 vccd1 vccd1 _14146_/CLK sky130_fd_sc_hd__buf_12
XFILLER_6_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08798_ _13666_/Q _08792_/X _08560_/X _08793_/X _08794_/X vssd1 vssd1 vccd1 vccd1
+ _13666_/D sky130_fd_sc_hd__o221a_1
Xrepeater682 _13370_/CLK vssd1 vssd1 vccd1 vccd1 _13368_/CLK sky130_fd_sc_hd__buf_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater693 _12635_/S vssd1 vssd1 vccd1 vccd1 _12610_/S sky130_fd_sc_hd__buf_8
XPHY_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ _08140_/A vssd1 vssd1 vccd1 vccd1 _07749_/X sky130_fd_sc_hd__buf_6
XPHY_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10760_ _10758_/Y _10691_/X _10759_/Y _10693_/X vssd1 vssd1 vccd1 vccd1 _10760_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09419_ _09419_/A _13023_/X vssd1 vssd1 vccd1 vccd1 _13318_/D sky130_fd_sc_hd__and2_1
XFILLER_164_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _11401_/A vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _12429_/X _06893_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12430_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12361_ _12360_/X _13202_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12361_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14100_ _14100_/CLK _14100_/D vssd1 vssd1 vccd1 vccd1 _14100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11312_ _11293_/X _11312_/B _11312_/C _11312_/D vssd1 vssd1 vccd1 vccd1 _11313_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12292_ _11699_/Y _14551_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12292_/X sky130_fd_sc_hd__mux2_2
XFILLER_49_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14031_ _14119_/CLK _14031_/D vssd1 vssd1 vccd1 vccd1 _14031_/Q sky130_fd_sc_hd__dfxtp_1
X_11243_ _14113_/Q vssd1 vssd1 vccd1 vccd1 _11243_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11174_ _14229_/Q _11170_/X _14424_/Q _11171_/X _11173_/X vssd1 vssd1 vccd1 vccd1
+ _11229_/B sky130_fd_sc_hd__a221oi_2
XFILLER_62_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10125_ _10125_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _12446_/S sky130_fd_sc_hd__or2_1
XFILLER_7_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10056_ _13358_/Q _09974_/B _09975_/A vssd1 vssd1 vccd1 vccd1 _10056_/X sky130_fd_sc_hd__o21a_1
XPHY_7473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13815_ _14130_/CLK _13815_/D vssd1 vssd1 vccd1 vccd1 _13815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13746_ _14121_/CLK _13746_/D vssd1 vssd1 vccd1 vccd1 _13746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10958_ _11430_/A vssd1 vssd1 vccd1 vccd1 _10958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13677_ _14146_/CLK _13677_/D vssd1 vssd1 vccd1 vccd1 _13677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10889_ _13950_/Q vssd1 vssd1 vccd1 vccd1 _10889_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12628_ _09839_/X _13330_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12628_/X sky130_fd_sc_hd__mux2_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12559_ _09953_/Y _13301_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12559_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14229_ _14495_/CLK _14229_/D vssd1 vssd1 vccd1 vccd1 _14229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09770_ _09770_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__or2_2
XFILLER_45_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06982_ _14566_/Q vssd1 vssd1 vccd1 vccd1 _06982_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08721_ _13709_/Q _08714_/X _08549_/X _08715_/X _08720_/X vssd1 vssd1 vccd1 vccd1
+ _13709_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _13745_/Q _08643_/X _08574_/X _08644_/X _08646_/X vssd1 vssd1 vccd1 vccd1
+ _13745_/D sky130_fd_sc_hd__o221a_1
X_07603_ _14263_/Q _07597_/X _07456_/X _07598_/X _07601_/X vssd1 vssd1 vccd1 vccd1
+ _14263_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08583_ _13780_/Q _08486_/A _08268_/X _08488_/A _08575_/X vssd1 vssd1 vccd1 vccd1
+ _13780_/D sky130_fd_sc_hd__o221a_1
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07534_ _14300_/Q _07532_/X _07374_/X _07533_/X _07527_/X vssd1 vssd1 vccd1 vccd1
+ _14300_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07465_ _14336_/Q _07459_/X _07381_/X _07460_/X _07461_/X vssd1 vssd1 vccd1 vccd1
+ _14336_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09204_ _09257_/A vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07396_ _08183_/A vssd1 vssd1 vccd1 vccd1 _07396_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _09135_/A vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ _09119_/A vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__buf_2
XFILLER_198_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08017_ _08017_/A vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__buf_2
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09968_ _13355_/Q _10052_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _13606_/Q _08916_/X _08917_/X _08918_/X _08910_/X vssd1 vssd1 vccd1 vccd1
+ _13606_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _09899_/A _09899_/B vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__or2_2
XPHY_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11930_ _14362_/Q vssd1 vssd1 vccd1 vccd1 _11930_/Y sky130_fd_sc_hd__inv_2
XPHY_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11861_ _13495_/Q vssd1 vssd1 vccd1 vccd1 _11861_/Y sky130_fd_sc_hd__inv_2
XPHY_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13600_ _14305_/CLK _13600_/D vssd1 vssd1 vccd1 vccd1 _13600_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _14104_/Q vssd1 vssd1 vccd1 vccd1 _10812_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14621_/CLK _14580_/D vssd1 vssd1 vccd1 vccd1 _14580_/Q sky130_fd_sc_hd__dfxtp_1
X_11792_ _13774_/Q vssd1 vssd1 vccd1 vccd1 _11792_/Y sky130_fd_sc_hd__inv_2
XPHY_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13531_ _14094_/CLK _13531_/D vssd1 vssd1 vccd1 vccd1 _13531_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _10734_/Y _10735_/X _10736_/Y _10737_/X _10742_/X vssd1 vssd1 vccd1 vccd1
+ _10754_/C sky130_fd_sc_hd__o221a_1
XFILLER_14_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ _14173_/CLK _13462_/D vssd1 vssd1 vccd1 vccd1 _13462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10674_ _14179_/Q vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12413_ _13216_/Q _06565_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12413_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13393_ _14183_/CLK _13393_/D vssd1 vssd1 vccd1 vccd1 _13393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ _13191_/Q _06853_/Y _12368_/S vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12275_ _12067_/Y _13376_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12275_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14014_ _14047_/CLK _14014_/D vssd1 vssd1 vccd1 vccd1 _14014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11226_ _11222_/Y _11223_/X _11224_/Y _11225_/X vssd1 vssd1 vccd1 vccd1 _11226_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11157_ _11152_/Y _10983_/X _11153_/Y _10985_/X _11156_/X vssd1 vssd1 vccd1 vccd1
+ _11158_/D sky130_fd_sc_hd__o221a_1
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10108_ _10138_/B _10143_/A vssd1 vssd1 vccd1 vccd1 _12467_/S sky130_fd_sc_hd__or2_1
XFILLER_49_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11088_ _13876_/Q vssd1 vssd1 vccd1 vccd1 _11088_/Y sky130_fd_sc_hd__inv_2
XPHY_7270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput260 la_oenb[69] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_hd__buf_1
XFILLER_62_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput271 la_oenb[79] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_hd__buf_1
XFILLER_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput282 la_oenb[89] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_hd__buf_1
X_10039_ _13360_/Q _09978_/B _09979_/A vssd1 vssd1 vccd1 vccd1 _10039_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput293 la_oenb[99] vssd1 vssd1 vccd1 vccd1 input293/X sky130_fd_sc_hd__buf_1
XFILLER_110_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13729_ _14056_/CLK _13729_/D vssd1 vssd1 vccd1 vccd1 _13729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ _07213_/A vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_203_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _09847_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _12888_/S sky130_fd_sc_hd__and2_2
XFILLER_138_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09753_ _13335_/Q vssd1 vssd1 vccd1 vccd1 _09785_/A sky130_fd_sc_hd__inv_2
XFILLER_210_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06965_ _06956_/X _12311_/X _06964_/Y _06958_/X vssd1 vssd1 vccd1 vccd1 _06966_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08704_ _08728_/A vssd1 vssd1 vccd1 vccd1 _08704_/X sky130_fd_sc_hd__buf_2
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _09684_/A vssd1 vssd1 vccd1 vccd1 _09684_/Y sky130_fd_sc_hd__inv_2
X_06896_ _14589_/Q vssd1 vssd1 vccd1 vccd1 _06897_/A sky130_fd_sc_hd__inv_2
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08635_ _08635_/A vssd1 vssd1 vccd1 vccd1 _08635_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08566_ input96/X vssd1 vssd1 vccd1 vccd1 _08566_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07517_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08497_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ _14346_/Q _07440_/X _07356_/X _07441_/X _07444_/X vssd1 vssd1 vccd1 vccd1
+ _14346_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07379_ _08167_/A vssd1 vssd1 vccd1 vccd1 _07379_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _13509_/Q _09111_/X _08967_/X _09112_/X _09117_/X vssd1 vssd1 vccd1 vccd1
+ _13509_/D sky130_fd_sc_hd__o221a_1
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _13940_/Q vssd1 vssd1 vccd1 vccd1 _10390_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09049_/A vssd1 vssd1 vccd1 vccd1 _09049_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _09789_/A _12057_/X _09901_/A _12058_/X vssd1 vssd1 vccd1 vccd1 _12060_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11011_ _11009_/Y _10952_/X _11010_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12962_ _12961_/X _12560_/X _12974_/S vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__mux2_1
XPHY_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11913_ _11908_/Y _10150_/A _11909_/Y _10153_/A _11912_/X vssd1 vssd1 vccd1 vccd1
+ _11948_/A sky130_fd_sc_hd__o221a_2
XPHY_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12534_/X _12892_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11834_/Y _11646_/X _11837_/X _11840_/X _11843_/X vssd1 vssd1 vccd1 vccd1
+ _11866_/C sky130_fd_sc_hd__o2111a_4
X_14632_ _14633_/CLK _14632_/D vssd1 vssd1 vccd1 vccd1 _14632_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14573_/CLK _14563_/D vssd1 vssd1 vccd1 vccd1 _14563_/Q sky130_fd_sc_hd__dfxtp_1
X_11775_ _13929_/Q vssd1 vssd1 vccd1 vccd1 _11775_/Y sky130_fd_sc_hd__inv_2
XPHY_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10726_ _14336_/Q vssd1 vssd1 vccd1 vccd1 _10726_/Y sky130_fd_sc_hd__inv_2
X_13514_ _14110_/CLK _13514_/D vssd1 vssd1 vccd1 vccd1 _13514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14494_ _14495_/CLK _14494_/D vssd1 vssd1 vccd1 vccd1 _14494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13445_ _14188_/CLK _13445_/D vssd1 vssd1 vccd1 vccd1 _13445_/Q sky130_fd_sc_hd__dfxtp_1
X_10657_ _13828_/Q vssd1 vssd1 vccd1 vccd1 _10657_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13376_ _14573_/CLK _13376_/D vssd1 vssd1 vccd1 vccd1 _13376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ _10586_/Y _10484_/X _10587_/Y _10487_/X vssd1 vssd1 vccd1 vccd1 _10588_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_122_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12327_ _13197_/Q _12326_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12258_ _12042_/Y _13359_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11209_ _11445_/A vssd1 vssd1 vccd1 vccd1 _11209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12189_ vssd1 vssd1 vccd1 vccd1 _12189_/HI _12189_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _14628_/Q _06733_/X _06748_/X _06726_/X _06749_/X vssd1 vssd1 vccd1 vccd1
+ _14628_/D sky130_fd_sc_hd__o221a_1
XFILLER_114_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06681_ _06679_/X _06680_/X _06679_/X _06680_/X vssd1 vssd1 vccd1 vccd1 _06682_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ _13855_/Q _08415_/X _08101_/X _08417_/X _08406_/X vssd1 vssd1 vccd1 vccd1
+ _13855_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _13893_/Q _08344_/X _08103_/X _08346_/X _08349_/X vssd1 vssd1 vccd1 vccd1
+ _13893_/D sky130_fd_sc_hd__o221a_1
XFILLER_204_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07302_ _14404_/Q _07238_/A _07083_/X _07240_/A _07301_/X vssd1 vssd1 vccd1 vccd1
+ _14404_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08282_ _13931_/Q _08274_/X _08105_/X _08276_/X _08278_/X vssd1 vssd1 vccd1 vccd1
+ _13931_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ _09063_/C vssd1 vssd1 vccd1 vccd1 _08744_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07164_ _07164_/A vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07095_ _14520_/Q _07092_/X _07015_/X _07094_/X _07079_/X vssd1 vssd1 vccd1 vccd1
+ _14520_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput520 _12149_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput531 _12159_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__clkbuf_2
Xoutput542 _12169_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput553 _12179_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput564 _12189_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__clkbuf_2
Xoutput575 _14639_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__clkbuf_2
XFILLER_132_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput586 _13274_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput597 _13284_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09805_ _09805_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__or2_2
XFILLER_64_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07997_ _14068_/Q _07991_/X _07852_/X _07992_/X _07995_/X vssd1 vssd1 vccd1 vccd1
+ _14068_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09736_ _10060_/A _12507_/S vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__nand2_1
X_06948_ _06954_/A _06948_/B vssd1 vssd1 vccd1 vccd1 _14576_/D sky130_fd_sc_hd__nor2_1
XFILLER_186_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09667_ _09657_/X _09666_/X _09657_/X _09666_/X vssd1 vssd1 vccd1 vccd1 _09667_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06879_ _09650_/A vssd1 vssd1 vccd1 vccd1 _06956_/A sky130_fd_sc_hd__buf_2
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08635_/A vssd1 vssd1 vccd1 vccd1 _08618_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09598_ _09557_/A _09597_/X _13255_/Q _09545_/A vssd1 vssd1 vccd1 vccd1 _13223_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08549_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__buf_4
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11560_ _13886_/Q vssd1 vssd1 vccd1 vccd1 _11560_/Y sky130_fd_sc_hd__inv_2
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10511_ _11693_/A vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__buf_6
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _14391_/Q vssd1 vssd1 vccd1 vccd1 _11491_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13352_/CLK _13230_/D vssd1 vssd1 vccd1 vccd1 _13262_/Q sky130_fd_sc_hd__dfxtp_2
X_10442_ _14214_/Q _10437_/X _14409_/Q _10438_/X _10441_/X vssd1 vssd1 vccd1 vccd1
+ _10519_/B sky130_fd_sc_hd__a221oi_2
XFILLER_87_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13161_ _12659_/X _13160_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__mux2_1
X_10373_ _10368_/Y _10228_/X _10369_/Y _10231_/X _10372_/X vssd1 vssd1 vccd1 vccd1
+ _10380_/C sky130_fd_sc_hd__o221a_1
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ vssd1 vssd1 vccd1 vccd1 _12112_/HI _12112_/LO sky130_fd_sc_hd__conb_1
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13092_ _12625_/X input334/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__buf_2
XFILLER_26_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _14110_/CLK _13994_/D vssd1 vssd1 vccd1 vccd1 _13994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12945_ _12553_/X _12944_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12945_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ _12530_/X input340/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12876_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_151 _11667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_162 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 input331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ _14627_/CLK _14615_/D vssd1 vssd1 vccd1 vccd1 _14615_/Q sky130_fd_sc_hd__dfxtp_1
X_11827_ _13651_/Q vssd1 vssd1 vccd1 vccd1 _11827_/Y sky130_fd_sc_hd__inv_2
XPHY_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 input337/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 input358/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11758_ _13532_/Q vssd1 vssd1 vccd1 vccd1 _11758_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14546_ _14611_/CLK _14546_/D vssd1 vssd1 vccd1 vccd1 _14546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ _11419_/A vssd1 vssd1 vccd1 vccd1 _10709_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14477_ _14481_/CLK _14477_/D vssd1 vssd1 vccd1 vccd1 _14477_/Q sky130_fd_sc_hd__dfxtp_1
X_11689_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__buf_2
XFILLER_31_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13428_ _14139_/CLK _13428_/D vssd1 vssd1 vccd1 vccd1 _13428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13359_ _14639_/CLK _13359_/D vssd1 vssd1 vccd1 vccd1 _13359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07920_ _14110_/Q _07918_/X _07759_/X _07919_/X _07913_/X vssd1 vssd1 vccd1 vccd1
+ _14110_/D sky130_fd_sc_hd__o221a_1
XFILLER_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07851_ _14147_/Q _07845_/X _07764_/X _07846_/X _07848_/X vssd1 vssd1 vccd1 vccd1
+ _14147_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06802_ _07130_/A vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__buf_4
XFILLER_211_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_07782_ _14179_/Q _07770_/X _07780_/X _07772_/X _07781_/X vssd1 vssd1 vccd1 vccd1
+ _14179_/D sky130_fd_sc_hd__o221a_1
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09521_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__clkbuf_2
X_06733_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06733_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09452_ _09456_/A _12935_/X vssd1 vssd1 vccd1 vccd1 _13292_/D sky130_fd_sc_hd__and2_1
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06664_ _06569_/Y _06663_/X _06569_/Y _06663_/X vssd1 vssd1 vccd1 vccd1 _06664_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _13862_/Q _08396_/X _08183_/X _08397_/X _08400_/X vssd1 vssd1 vccd1 vccd1
+ _13862_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__buf_2
XFILLER_209_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06595_ _06595_/A vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__clkbuf_4
X_08334_ _13900_/Q _08274_/A _08186_/X _08276_/A _08329_/X vssd1 vssd1 vccd1 vccd1
+ _13900_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08265_ _13939_/Q _08198_/A _08186_/X _08201_/A _08264_/X vssd1 vssd1 vccd1 vccd1
+ _13939_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07216_ _14452_/Q _07209_/X _06820_/X _07210_/X _07213_/X vssd1 vssd1 vccd1 vccd1
+ _14452_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08196_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__inv_2
XFILLER_179_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07147_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07147_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07078_ _07130_/A vssd1 vssd1 vccd1 vccd1 _07122_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput372 _12209_/X vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput383 _12219_/X vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput394 _12229_/X vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09719_ _14581_/Q _06933_/Y _06927_/Y _14579_/Q vssd1 vssd1 vccd1 vccd1 _09719_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10991_ _10982_/Y _10983_/X _10984_/Y _10985_/X _10990_/X vssd1 vssd1 vccd1 vccd1
+ _10992_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _09578_/X _12729_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _13346_/Q _12660_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14400_ _14633_/CLK _14400_/D vssd1 vssd1 vccd1 vccd1 _14400_/Q sky130_fd_sc_hd__dfxtp_1
X_11612_ _14511_/Q vssd1 vssd1 vccd1 vccd1 _11612_/Y sky130_fd_sc_hd__inv_2
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _13317_/Q _12591_/X _12655_/S vssd1 vssd1 vccd1 vccd1 _12592_/X sky130_fd_sc_hd__mux2_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ _14527_/CLK _14331_/D vssd1 vssd1 vccd1 vccd1 _14331_/Q sky130_fd_sc_hd__dfxtp_1
X_11543_ _14158_/Q vssd1 vssd1 vccd1 vccd1 _11543_/Y sky130_fd_sc_hd__inv_2
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14305_/CLK _14262_/D vssd1 vssd1 vccd1 vccd1 _14262_/Q sky130_fd_sc_hd__dfxtp_1
X_11474_ _13962_/Q vssd1 vssd1 vccd1 vccd1 _11474_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13213_ _14459_/CLK _13213_/D vssd1 vssd1 vccd1 vccd1 _13213_/Q sky130_fd_sc_hd__dfxtp_4
X_10425_ _11397_/A vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _14305_/CLK _14193_/D vssd1 vssd1 vccd1 vccd1 _14193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ _12651_/X input337/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__mux2_1
X_10356_ _13978_/Q vssd1 vssd1 vccd1 vccd1 _10356_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13075_ _12616_/X _13074_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10287_ _14171_/Q vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12026_ _14481_/Q vssd1 vssd1 vccd1 vccd1 _12026_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13977_ _14095_/CLK _13977_/D vssd1 vssd1 vccd1 vccd1 _13977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12928_ _12545_/X input358/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12525_/X _12858_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14529_ _14529_/CLK _14529_/D vssd1 vssd1 vccd1 vccd1 _14529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08050_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__buf_2
XFILLER_204_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07001_ _07004_/A _07001_/B vssd1 vssd1 vccd1 vccd1 _14561_/D sky130_fd_sc_hd__nor2_1
XFILLER_122_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08952_ _13594_/Q _08944_/X _08950_/X _08946_/X _08951_/X vssd1 vssd1 vccd1 vccd1
+ _13594_/D sky130_fd_sc_hd__o221a_1
XFILLER_48_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07903_ _07927_/A vssd1 vssd1 vccd1 vccd1 _07903_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08883_ _13622_/Q _08876_/X _08572_/X _08877_/X _08880_/X vssd1 vssd1 vccd1 vccd1
+ _13622_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07834_ _14157_/Q _07829_/X _07738_/X _07830_/X _07831_/X vssd1 vssd1 vccd1 vccd1
+ _14157_/D sky130_fd_sc_hd__o221a_1
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07765_ _14186_/Q _07758_/X _07764_/X _07760_/X _07756_/X vssd1 vssd1 vccd1 vccd1
+ _14186_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06716_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06716_/X sky130_fd_sc_hd__clkbuf_2
X_09504_ _13259_/Q _09500_/X _12254_/X _09501_/X vssd1 vssd1 vccd1 vccd1 _13259_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07696_ _14211_/Q _07634_/A _07401_/X _07636_/A _07692_/X vssd1 vssd1 vccd1 vccd1
+ _14211_/D sky130_fd_sc_hd__o221a_1
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09435_ _09438_/A _13007_/X vssd1 vssd1 vccd1 vccd1 _13306_/D sky130_fd_sc_hd__and2_1
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06647_ _06626_/A _06561_/A _06625_/Y _06561_/Y vssd1 vssd1 vccd1 vccd1 _06647_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09366_ _09370_/A _12847_/X vssd1 vssd1 vccd1 vccd1 _13362_/D sky130_fd_sc_hd__and2_1
XFILLER_55_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06578_ _06574_/Y _06575_/Y _08977_/A _08983_/A vssd1 vssd1 vccd1 vccd1 _06578_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08317_ _13911_/Q _08310_/X _08158_/X _08311_/X _08313_/X vssd1 vssd1 vccd1 vccd1
+ _13911_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_40 _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _13410_/Q _09294_/X _08126_/A _09295_/X _09290_/X vssd1 vssd1 vccd1 vccd1
+ _13410_/D sky130_fd_sc_hd__o221a_1
XFILLER_166_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_51 _07759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 _07825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08248_ _08383_/A vssd1 vssd1 vccd1 vccd1 _08288_/A sky130_fd_sc_hd__buf_6
XANTENNA_73 _08167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_84 _08558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_95 _08942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08179_ _08179_/A vssd1 vssd1 vccd1 vccd1 _08179_/X sky130_fd_sc_hd__buf_4
XFILLER_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10210_ _13539_/Q _10206_/X _13780_/Q _10209_/X vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11190_ _11426_/A vssd1 vssd1 vccd1 vccd1 _11190_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10141_ _10141_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _12425_/S sky130_fd_sc_hd__or2_1
XFILLER_0_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10072_ _10079_/A _10118_/A vssd1 vssd1 vccd1 vccd1 _12497_/S sky130_fd_sc_hd__or2_1
XFILLER_118_1884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13900_ _14169_/CLK _13900_/D vssd1 vssd1 vccd1 vccd1 _13900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13831_ _14107_/CLK _13831_/D vssd1 vssd1 vccd1 vccd1 _13831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13762_ _13996_/CLK _13762_/D vssd1 vssd1 vccd1 vccd1 _13762_/Q sky130_fd_sc_hd__dfxtp_1
X_10974_ _13593_/Q vssd1 vssd1 vccd1 vccd1 _10974_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ _09567_/X _12712_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12713_/X sky130_fd_sc_hd__mux2_1
X_13693_ _14056_/CLK _13693_/D vssd1 vssd1 vccd1 vccd1 _13693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _09826_/X _13338_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__mux2_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _09941_/Y _13309_/Q _12603_/S vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314_ _14527_/CLK _14314_/D vssd1 vssd1 vccd1 vccd1 _14314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ _11524_/Y _11424_/X _11525_/Y _11426_/X vssd1 vssd1 vccd1 vccd1 _11526_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14245_ _14325_/CLK _14245_/D vssd1 vssd1 vccd1 vccd1 _14245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _11457_/A vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10408_ _10403_/Y _10214_/X _10404_/Y _10217_/X _10407_/X vssd1 vssd1 vccd1 vccd1
+ _10421_/B sky130_fd_sc_hd__o221a_4
X_14176_ _14178_/CLK _14176_/D vssd1 vssd1 vccd1 vccd1 _14176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ _13921_/Q vssd1 vssd1 vccd1 vccd1 _11388_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10339_ _10320_/X _10339_/B _10339_/C _10339_/D vssd1 vssd1 vccd1 vccd1 _10340_/D
+ sky130_fd_sc_hd__and4b_1
X_13127_ _12641_/X _13126_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13058_ _13057_/X _12608_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12009_ _13577_/Q _10206_/A _13818_/Q _10209_/A vssd1 vssd1 vccd1 vccd1 _12009_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07550_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07550_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06501_ _06512_/A _06509_/C vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__or2_1
XFILLER_207_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07481_ _14326_/Q _07411_/A _07480_/X _07414_/A _07476_/X vssd1 vssd1 vccd1 vccd1
+ _14326_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _13454_/Q _09215_/X _07723_/A _09217_/X _09219_/X vssd1 vssd1 vccd1 vccd1
+ _13454_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09151_ _13493_/Q _09146_/X _08837_/X _09148_/X _09149_/X vssd1 vssd1 vccd1 vccd1
+ _13493_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08102_ _14011_/Q _08095_/X _08101_/X _08097_/X _08089_/X vssd1 vssd1 vccd1 vccd1
+ _14011_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09082_ _13531_/Q _09077_/X _09009_/X _09079_/X _09074_/X vssd1 vssd1 vccd1 vccd1
+ _13531_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08033_ _14049_/Q _08025_/X _07712_/X _08027_/X _08032_/X vssd1 vssd1 vccd1 vccd1
+ _14049_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput60 la_data_in[119] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_1
Xinput71 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_1
XFILLER_200_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput82 la_data_in[23] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_1
XFILLER_11_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput93 la_data_in[33] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09984_ _13363_/Q _09984_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08935_ _08935_/A vssd1 vssd1 vccd1 vccd1 _08935_/X sky130_fd_sc_hd__buf_6
XFILLER_83_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08866_ _13632_/Q _08860_/X _08632_/X _08861_/X _08863_/X vssd1 vssd1 vccd1 vccd1
+ _13632_/D sky130_fd_sc_hd__o221a_1
XPHY_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater650 _14529_/CLK vssd1 vssd1 vccd1 vccd1 _14527_/CLK sky130_fd_sc_hd__buf_12
XPHY_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07817_ _14165_/Q _07808_/X _07714_/X _07811_/X _07812_/X vssd1 vssd1 vccd1 vccd1
+ _14165_/D sky130_fd_sc_hd__o221a_1
Xrepeater661 _14095_/CLK vssd1 vssd1 vccd1 vccd1 _14100_/CLK sky130_fd_sc_hd__buf_8
XFILLER_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _13667_/Q _08792_/X _08558_/X _08793_/X _08794_/X vssd1 vssd1 vccd1 vccd1
+ _13667_/D sky130_fd_sc_hd__o221a_1
Xrepeater672 _14071_/CLK vssd1 vssd1 vccd1 vccd1 _14143_/CLK sky130_fd_sc_hd__buf_12
Xrepeater683 _12231_/A vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__buf_12
XPHY_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater694 input39/X vssd1 vssd1 vccd1 vccd1 _12635_/S sky130_fd_sc_hd__buf_8
XFILLER_211_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07748_ _14193_/Q _07745_/X _07746_/X _07747_/X _07743_/X vssd1 vssd1 vccd1 vccd1
+ _14193_/D sky130_fd_sc_hd__o221a_1
XFILLER_183_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07679_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07679_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09418_ _09419_/A _13083_/X vssd1 vssd1 vccd1 vccd1 _13319_/D sky130_fd_sc_hd__and2_1
X_10690_ _13666_/Q vssd1 vssd1 vccd1 vccd1 _10690_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09349_ _09351_/A _12923_/X vssd1 vssd1 vccd1 vccd1 _13375_/D sky130_fd_sc_hd__and2_1
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12360_ _13202_/Q _12359_/X input78/X vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _11306_/Y _11219_/X _11307_/Y _11221_/X _11310_/X vssd1 vssd1 vccd1 vccd1
+ _11312_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12291_ _11740_/Y _14552_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__mux2_2
XFILLER_120_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14030_ _14119_/CLK _14030_/D vssd1 vssd1 vccd1 vccd1 _14030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11242_ _13840_/Q vssd1 vssd1 vccd1 vccd1 _11242_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _13403_/Q _11042_/X _13715_/Q _11172_/X vssd1 vssd1 vccd1 vccd1 _11173_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_84_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10124_ _10138_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__buf_1
XFILLER_27_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ _13357_/Q _09972_/B _09973_/A vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__o21a_1
XPHY_7463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ _14130_/CLK _13814_/D vssd1 vssd1 vccd1 vccd1 _13814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13745_ _14094_/CLK _13745_/D vssd1 vssd1 vccd1 vccd1 _13745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10957_ _11429_/A vssd1 vssd1 vccd1 vccd1 _10957_/X sky130_fd_sc_hd__buf_2
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13676_ _14146_/CLK _13676_/D vssd1 vssd1 vccd1 vccd1 _13676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10888_ _14223_/Q _10696_/X _14418_/Q _10697_/X _10887_/X vssd1 vssd1 vccd1 vccd1
+ _10921_/B sky130_fd_sc_hd__a221oi_2
XFILLER_164_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12627_ _13331_/Q _12626_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12627_/X sky130_fd_sc_hd__mux2_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12558_ _13302_/Q _12557_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12558_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _13449_/Q vssd1 vssd1 vccd1 vccd1 _11509_/Y sky130_fd_sc_hd__inv_2
X_12489_ _12488_/X _06970_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12489_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14228_ _14495_/CLK _14228_/D vssd1 vssd1 vccd1 vccd1 _14228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14470_/CLK _14159_/D vssd1 vssd1 vccd1 vccd1 _14159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06981_ _06991_/A _06981_/B vssd1 vssd1 vccd1 vccd1 _14567_/D sky130_fd_sc_hd__nor2_1
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08720_ _08728_/A vssd1 vssd1 vccd1 vccd1 _08720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08651_ _13746_/Q _08643_/X _08572_/X _08644_/X _08646_/X vssd1 vssd1 vccd1 vccd1
+ _13746_/D sky130_fd_sc_hd__o221a_1
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07602_ _14264_/Q _07597_/X _07367_/X _07598_/X _07601_/X vssd1 vssd1 vccd1 vccd1
+ _14264_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08582_ _13781_/Q _08486_/A _08581_/X _08488_/A _08575_/X vssd1 vssd1 vccd1 vccd1
+ _13781_/D sky130_fd_sc_hd__o221a_1
XFILLER_19_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07533_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07533_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07464_ _14337_/Q _07459_/X _07379_/X _07460_/X _07461_/X vssd1 vssd1 vccd1 vccd1
+ _14337_/D sky130_fd_sc_hd__o221a_1
XFILLER_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09203_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__inv_2
XFILLER_91_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07395_ _14370_/Q _07387_/X _07394_/X _07389_/X _07385_/X vssd1 vssd1 vccd1 vccd1
+ _14370_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09134_ _09188_/A vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09065_ _09120_/A vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__inv_2
XFILLER_190_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08016_ _14055_/Q _07955_/A _07798_/X _07957_/A _08011_/X vssd1 vssd1 vccd1 vccd1
+ _14055_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _13353_/Q _09967_/B _13354_/Q vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__and3_1
XFILLER_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08918_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09898_ _09898_/A _09931_/A vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__or2_2
XPHY_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _13643_/Q _08844_/X _08519_/X _08845_/X _08847_/X vssd1 vssd1 vccd1 vccd1
+ _13643_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11860_ _14165_/Q vssd1 vssd1 vccd1 vccd1 _11860_/Y sky130_fd_sc_hd__inv_2
XPHY_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _13831_/Q vssd1 vssd1 vccd1 vccd1 _10811_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11791_ _13969_/Q vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__inv_2
XPHY_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13530_ _14094_/CLK _13530_/D vssd1 vssd1 vccd1 vccd1 _13530_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _10738_/Y _10739_/X _10740_/Y _10741_/X vssd1 vssd1 vccd1 vccd1 _10742_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ _14173_/CLK _13461_/D vssd1 vssd1 vccd1 vccd1 _13461_/Q sky130_fd_sc_hd__dfxtp_1
X_10673_ _13587_/Q vssd1 vssd1 vccd1 vccd1 _10673_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12412_ _12411_/X _13217_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13392_ _14183_/CLK _13392_/D vssd1 vssd1 vccd1 vccd1 _13392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343_ _12342_/X _13192_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ _12066_/Y _13375_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12274_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ _14130_/CLK _14013_/D vssd1 vssd1 vccd1 vccd1 _14013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11225_ _11461_/A vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11156_ _11154_/Y _10987_/X _11155_/Y _10989_/X vssd1 vssd1 vccd1 vccd1 _11156_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__or2_1
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11087_ _13759_/Q vssd1 vssd1 vccd1 vccd1 _11087_/Y sky130_fd_sc_hd__inv_2
XPHY_7260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput250 la_oenb[5] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__buf_1
XFILLER_209_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput261 la_oenb[6] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_hd__buf_1
XPHY_7282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput272 la_oenb[7] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_hd__buf_1
X_10038_ _13359_/Q _09976_/B _09977_/A vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__o21a_1
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput283 la_oenb[8] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_1
XFILLER_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput294 la_oenb[9] vssd1 vssd1 vccd1 vccd1 input294/X sky130_fd_sc_hd__buf_1
XFILLER_64_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11989_ _11989_/A _11989_/B _11989_/C _11989_/D vssd1 vssd1 vccd1 vccd1 _11989_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_166_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _14047_/CLK _13728_/D vssd1 vssd1 vccd1 vccd1 _13728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13659_ _14047_/CLK _13659_/D vssd1 vssd1 vccd1 vccd1 _13659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07180_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09821_ _09785_/A _09785_/B _09820_/Y vssd1 vssd1 vccd1 vccd1 _09821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09752_ _13336_/Q vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__inv_2
X_06964_ _14571_/Q vssd1 vssd1 vccd1 vccd1 _06964_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08703_ _13720_/Q _08698_/X _08521_/X _08699_/X _08696_/X vssd1 vssd1 vccd1 vccd1
+ _13720_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09683_ _06952_/Y _14572_/Q _14574_/Q _06961_/Y vssd1 vssd1 vccd1 vccd1 _09684_/A
+ sky130_fd_sc_hd__o22a_1
X_06895_ _06899_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _14590_/D sky130_fd_sc_hd__nor2_1
XFILLER_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08634_ _13755_/Q _08626_/X _08549_/X _08627_/X _08628_/X vssd1 vssd1 vccd1 vccd1
+ _13755_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08565_/A vssd1 vssd1 vccd1 vccd1 _08565_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07516_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07516_/X sky130_fd_sc_hd__clkbuf_2
X_08496_ _08829_/A vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__buf_2
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07447_ _14347_/Q _07440_/X _07354_/X _07441_/X _07444_/X vssd1 vssd1 vccd1 vccd1
+ _14347_/D sky130_fd_sc_hd__o221a_1
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07378_ _14377_/Q _07373_/X _07377_/X _07375_/X _07371_/X vssd1 vssd1 vccd1 vccd1
+ _14377_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _09048_/A vssd1 vssd1 vccd1 vccd1 _09048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11010_ _13516_/Q vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12961_ _12560_/X _12960_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11912_ _11910_/Y _10156_/A _11911_/Y _10159_/A vssd1 vssd1 vccd1 vccd1 _11912_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12534_/X input354/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14631_ _14633_/CLK _14631_/D vssd1 vssd1 vccd1 vccd1 _14631_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11843_ _11841_/Y _11658_/X _11842_/Y _11660_/X vssd1 vssd1 vccd1 vccd1 _11843_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14573_/CLK _14562_/D vssd1 vssd1 vccd1 vccd1 _14562_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11774_ _11769_/Y _11679_/X _11770_/Y _11681_/X _11773_/X vssd1 vssd1 vccd1 vccd1
+ _11781_/C sky130_fd_sc_hd__o221a_1
XPHY_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _14110_/CLK _13513_/D vssd1 vssd1 vccd1 vccd1 _13513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10725_ _11435_/A vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__buf_2
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14493_ _14495_/CLK _14493_/D vssd1 vssd1 vccd1 vccd1 _14493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13444_ _14459_/CLK _13444_/D vssd1 vssd1 vccd1 vccd1 _13444_/Q sky130_fd_sc_hd__dfxtp_1
X_10656_ _10654_/Y _10448_/X _10655_/Y _10451_/X vssd1 vssd1 vccd1 vccd1 _10656_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10587_ _14372_/Q vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__inv_2
X_13375_ _14573_/CLK _13375_/D vssd1 vssd1 vccd1 vccd1 _13375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12326_ _13197_/Q input95/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12257_ _12041_/Y _13358_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12257_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _14307_/Q vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__inv_2
X_12188_ vssd1 vssd1 vccd1 vccd1 _12188_/HI _12188_/LO sky130_fd_sc_hd__conb_1
XFILLER_155_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11139_ _13210_/Q _11013_/X _14033_/Q _10957_/X _11138_/X vssd1 vssd1 vccd1 vccd1
+ _11139_/X sky130_fd_sc_hd__a221o_4
XFILLER_211_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06680_ input96/X _08974_/A _06637_/Y _06589_/Y vssd1 vssd1 vccd1 vccd1 _06680_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08350_ _13894_/Q _08344_/X _08101_/X _08346_/X _08349_/X vssd1 vssd1 vccd1 vccd1
+ _13894_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07301_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07301_/X sky130_fd_sc_hd__buf_2
XFILLER_149_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08281_ _13932_/Q _08274_/X _08103_/X _08276_/X _08278_/X vssd1 vssd1 vccd1 vccd1
+ _13932_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07232_ _07232_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _09063_/C sky130_fd_sc_hd__or2_2
XFILLER_14_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07163_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07164_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _07094_/A vssd1 vssd1 vccd1 vccd1 _07094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput510 _12140_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput521 _12150_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__clkbuf_2
Xoutput532 _12160_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput543 _12170_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__clkbuf_2
Xoutput554 _12180_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput565 _12190_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput576 _13255_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput587 _13256_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput598 _13257_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09804_ _13346_/Q vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__inv_2
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07996_ _14069_/Q _07991_/X _07764_/X _07992_/X _07995_/X vssd1 vssd1 vccd1 vccd1
+ _14069_/D sky130_fd_sc_hd__o221a_1
X_09735_ _12510_/S _10077_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06947_ _06937_/X _12306_/X _06946_/Y _06939_/X vssd1 vssd1 vccd1 vccd1 _06948_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09666_ _06912_/Y _14577_/Q _14585_/Q _06943_/A vssd1 vssd1 vccd1 vccd1 _09666_/X
+ sky130_fd_sc_hd__o22a_1
X_06878_ _06918_/A vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08617_ _13765_/Q _08610_/X _08523_/X _08611_/X _08612_/X vssd1 vssd1 vccd1 vccd1
+ _13765_/D sky130_fd_sc_hd__o221a_1
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09597_ _09597_/A _12346_/X vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__and2_1
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _13795_/Q _08540_/X _08243_/X _08542_/X _08538_/X vssd1 vssd1 vccd1 vccd1
+ _13795_/D sky130_fd_sc_hd__o221a_1
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08479_ _13820_/Q _08415_/A _08190_/X _08417_/A _08474_/X vssd1 vssd1 vccd1 vccd1
+ _13820_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10510_ _13466_/Q vssd1 vssd1 vccd1 vccd1 _10510_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _14625_/Q vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__inv_2
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10441_ _13388_/Q _10305_/X _13700_/Q _10440_/X vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _10370_/Y _10234_/X _10371_/Y _10237_/X vssd1 vssd1 vccd1 vccd1 _10372_/X
+ sky130_fd_sc_hd__o22a_1
X_13160_ _12659_/X input350/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13160_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12111_ vssd1 vssd1 vccd1 vccd1 _12111_/HI _12111_/LO sky130_fd_sc_hd__conb_1
X_13091_ _12623_/X _13090_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12042_ _09777_/A _12035_/X _09889_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12042_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13993_ _14107_/CLK _13993_/D vssd1 vssd1 vccd1 vccd1 _13993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12944_ _12553_/X input352/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12944_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12529_/X _12874_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_130 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_141 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_152 _11762_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14614_ _14627_/CLK _14614_/D vssd1 vssd1 vccd1 vccd1 _14614_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_163 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _13690_/Q vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 input331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_185 input341/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_196 input358/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14545_ _14611_/CLK _14545_/D vssd1 vssd1 vccd1 vccd1 _14545_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _14007_/Q vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _13829_/Q vssd1 vssd1 vccd1 vccd1 _10708_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14476_ _14481_/CLK _14476_/D vssd1 vssd1 vccd1 vccd1 _14476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11688_ _13927_/Q vssd1 vssd1 vccd1 vccd1 _11688_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13427_ _14139_/CLK _13427_/D vssd1 vssd1 vccd1 vccd1 _13427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10639_ _13469_/Q vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13358_ _14639_/CLK _13358_/D vssd1 vssd1 vccd1 vccd1 _13358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12309_ _10880_/Y _14534_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12309_/X sky130_fd_sc_hd__mux2_2
XFILLER_143_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13289_ _13996_/CLK _13289_/D vssd1 vssd1 vccd1 vccd1 _13289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07850_ _14148_/Q _07845_/X _07762_/X _07846_/X _07848_/X vssd1 vssd1 vccd1 vccd1
+ _14148_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06801_ _08158_/A vssd1 vssd1 vccd1 vccd1 _06801_/X sky130_fd_sc_hd__buf_4
XFILLER_81_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07781_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07781_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_133_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _09514_/X _09519_/X _13285_/Q _09517_/X vssd1 vssd1 vccd1 vccd1 _13253_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06732_ _06823_/A vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__buf_2
XFILLER_168_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06663_ _06639_/Y _08935_/A _08930_/A _06596_/Y vssd1 vssd1 vccd1 vccd1 _06663_/X
+ sky130_fd_sc_hd__o22a_1
X_09451_ _09451_/A vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08402_ _13863_/Q _08396_/X _08181_/X _08397_/X _08400_/X vssd1 vssd1 vccd1 vccd1
+ _13863_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09382_ _09382_/A _13159_/X vssd1 vssd1 vccd1 vccd1 _13348_/D sky130_fd_sc_hd__and2_1
X_06594_ _06596_/A vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08333_ _13901_/Q _08326_/X _08183_/X _08327_/X _08329_/X vssd1 vssd1 vccd1 vccd1
+ _13901_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08264_ _08288_/A vssd1 vssd1 vccd1 vccd1 _08264_/X sky130_fd_sc_hd__buf_4
XFILLER_18_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07215_ _14453_/Q _07209_/X _06817_/X _07210_/X _07213_/X vssd1 vssd1 vccd1 vccd1
+ _14453_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08195_ _08341_/A _11646_/A vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__or2_4
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07146_ _14490_/Q _07144_/X _06825_/X _07145_/X _07139_/X vssd1 vssd1 vccd1 vccd1
+ _14490_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07077_ _14525_/Q _07069_/X _06837_/X _07070_/X _07071_/X vssd1 vssd1 vccd1 vccd1
+ _14525_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput373 _12210_/X vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput384 _12220_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput395 _12230_/X vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07979_ _14079_/Q _07974_/X _07738_/X _07975_/X _07978_/X vssd1 vssd1 vccd1 vccd1
+ _14079_/D sky130_fd_sc_hd__o221a_1
XFILLER_169_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09718_ _06893_/X _09706_/X _06893_/A _09706_/X vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10990_ _10986_/Y _10987_/X _10988_/Y _10989_/X vssd1 vssd1 vccd1 vccd1 _10990_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _09620_/X _09648_/X _09620_/X _09648_/X vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_71_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _09806_/X _13346_/Q _12666_/S vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__mux2_1
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11611_ _13220_/Q _11485_/X _14043_/Q _11429_/X _11610_/X vssd1 vssd1 vccd1 vccd1
+ _11611_/X sky130_fd_sc_hd__a221o_4
XFILLER_19_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _09928_/Y _13317_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__mux2_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14330_ _14633_/CLK _14330_/D vssd1 vssd1 vccd1 vccd1 _14330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _13924_/Q vssd1 vssd1 vccd1 vccd1 _11542_/Y sky130_fd_sc_hd__inv_2
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14261_ _14305_/CLK _14261_/D vssd1 vssd1 vccd1 vccd1 _14261_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _14235_/Q _11406_/X _14430_/Q _11407_/X _11472_/X vssd1 vssd1 vccd1 vccd1
+ _11507_/B sky130_fd_sc_hd__a221oi_2
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13212_ _13370_/CLK _13212_/D vssd1 vssd1 vccd1 vccd1 _13212_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10424_ _11633_/A vssd1 vssd1 vccd1 vccd1 _11397_/A sky130_fd_sc_hd__buf_4
XFILLER_197_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14192_ _14305_/CLK _14192_/D vssd1 vssd1 vccd1 vccd1 _14192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13143_ _12649_/X _13142_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13143_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10355_ _10353_/Y _10188_/X _10354_/Y _10191_/X vssd1 vssd1 vccd1 vccd1 _10355_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10286_ _13579_/Q vssd1 vssd1 vccd1 vccd1 _10286_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13074_ _13073_/X _12616_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12025_ _13499_/Q vssd1 vssd1 vccd1 vccd1 _12025_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13976_ _14095_/CLK _13976_/D vssd1 vssd1 vccd1 vccd1 _13976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12927_ _12543_/X _12926_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12927_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12858_ _12525_/X _12857_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12858_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ _11804_/Y _11669_/X _11805_/Y _11671_/X _11808_/X vssd1 vssd1 vccd1 vccd1
+ _11822_/B sky130_fd_sc_hd__o221a_2
XFILLER_15_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ _09533_/X _12788_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12789_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14528_ _14529_/CLK _14528_/D vssd1 vssd1 vccd1 vccd1 _14528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14459_ _14459_/CLK _14459_/D vssd1 vssd1 vccd1 vccd1 _14459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07000_ _06857_/A _12321_/X _06999_/Y _06861_/A vssd1 vssd1 vccd1 vccd1 _07001_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08951_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07902_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08882_ _13623_/Q _08876_/X _08570_/X _08877_/X _08880_/X vssd1 vssd1 vccd1 vccd1
+ _13623_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07833_ _14158_/Q _07829_/X _07736_/X _07830_/X _07831_/X vssd1 vssd1 vccd1 vccd1
+ _14158_/D sky130_fd_sc_hd__o221a_1
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07764_ _08155_/A vssd1 vssd1 vccd1 vccd1 _07764_/X sky130_fd_sc_hd__buf_4
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _13260_/Q _09500_/X _12255_/X _09501_/X vssd1 vssd1 vccd1 vccd1 _13260_/D
+ sky130_fd_sc_hd__o22a_1
X_06715_ _06811_/A vssd1 vssd1 vccd1 vccd1 _06790_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07695_ _14212_/Q _07634_/A _07399_/X _07636_/A _07692_/X vssd1 vssd1 vccd1 vccd1
+ _14212_/D sky130_fd_sc_hd__o221a_1
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09434_ _09438_/A _13003_/X vssd1 vssd1 vccd1 vccd1 _13307_/D sky130_fd_sc_hd__and2_1
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06646_ _06553_/Y _06668_/A _08917_/A _06645_/Y vssd1 vssd1 vccd1 vccd1 _06646_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09365_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06577_ input92/X vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__buf_4
XFILLER_205_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08316_ _13912_/Q _08310_/X _08243_/X _08311_/X _08313_/X vssd1 vssd1 vccd1 vccd1
+ _13912_/D sky130_fd_sc_hd__o221a_1
X_09296_ _13411_/Q _09294_/X _08123_/A _09295_/X _09290_/X vssd1 vssd1 vccd1 vccd1
+ _13411_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_30 _06793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_41 _07362_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _07762_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_63 _07886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08247_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08247_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_74 _08169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_85 _08558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_96 _08948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08178_ _13982_/Q _08174_/X _07867_/X _08176_/X _08172_/X vssd1 vssd1 vccd1 vccd1
+ _13982_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07129_ _14500_/Q _07127_/X _06789_/X _07128_/X _07122_/X vssd1 vssd1 vccd1 vccd1
+ _14500_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10140_ _10140_/A _12509_/S vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10071_ _10113_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__or2_1
XFILLER_62_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13830_ _14107_/CLK _13830_/D vssd1 vssd1 vccd1 vccd1 _13830_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13761_ _13996_/CLK _13761_/D vssd1 vssd1 vccd1 vccd1 _13761_/Q sky130_fd_sc_hd__dfxtp_1
X_10973_ _11445_/A vssd1 vssd1 vccd1 vccd1 _10973_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _09567_/X input333/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__mux2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13692_ _14056_/CLK _13692_/D vssd1 vssd1 vccd1 vccd1 _13692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12643_ _13339_/Q _12642_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__mux2_1
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _13310_/Q _12573_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__mux2_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _14527_/CLK _14313_/D vssd1 vssd1 vccd1 vccd1 _14313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11525_ _13527_/Q vssd1 vssd1 vccd1 vccd1 _11525_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14244_ _14325_/CLK _14244_/D vssd1 vssd1 vccd1 vccd1 _14244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ _14156_/Q vssd1 vssd1 vccd1 vccd1 _11456_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10407_ _10405_/Y _10220_/X _10406_/Y _10223_/X vssd1 vssd1 vccd1 vccd1 _10407_/X
+ sky130_fd_sc_hd__o22a_1
X_14175_ _14178_/CLK _14175_/D vssd1 vssd1 vccd1 vccd1 _14175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11387_ _11382_/Y _11209_/X _11383_/Y _11211_/X _11386_/X vssd1 vssd1 vccd1 vccd1
+ _11394_/C sky130_fd_sc_hd__o221a_1
XFILLER_140_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13126_ _13125_/X _12641_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10338_ _10333_/Y _10242_/X _10334_/Y _10245_/X _10337_/X vssd1 vssd1 vccd1 vccd1
+ _10339_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13057_ _12608_/X _13056_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__mux2_1
X_10269_ _14093_/Q vssd1 vssd1 vccd1 vccd1 _10269_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12008_ _11998_/Y _10178_/A _12001_/X _12004_/X _12007_/X vssd1 vssd1 vccd1 vccd1
+ _12030_/C sky130_fd_sc_hd__o2111a_4
XFILLER_152_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13959_ _13996_/CLK _13959_/D vssd1 vssd1 vccd1 vccd1 _13959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06500_ _06500_/A _06510_/A vssd1 vssd1 vccd1 vccd1 _06509_/C sky130_fd_sc_hd__or2_1
X_07480_ _08268_/A vssd1 vssd1 vccd1 vccd1 _07480_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_185_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09150_ _13494_/Q _09146_/X _08833_/X _09148_/X _09149_/X vssd1 vssd1 vccd1 vccd1
+ _13494_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08101_ _08825_/A vssd1 vssd1 vccd1 vccd1 _08101_/X sky130_fd_sc_hd__buf_4
XFILLER_147_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09081_ _13532_/Q _09077_/X _08837_/X _09079_/X _09074_/X vssd1 vssd1 vccd1 vccd1
+ _13532_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08032_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08032_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_1
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_1
Xinput72 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_1
XFILLER_11_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput83 la_data_in[24] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_1
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput94 la_data_in[34] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_2
XFILLER_192_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _09983_/A vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__inv_2
XFILLER_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08934_ _13600_/Q _08929_/X _08933_/X _08931_/X _08923_/X vssd1 vssd1 vccd1 vccd1
+ _13600_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _13633_/Q _08860_/X _08546_/X _08861_/X _08863_/X vssd1 vssd1 vccd1 vccd1
+ _13633_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater640 _14459_/CLK vssd1 vssd1 vccd1 vccd1 _14538_/CLK sky130_fd_sc_hd__buf_12
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07816_ _14166_/Q _07808_/X _07712_/X _07811_/X _07812_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/D sky130_fd_sc_hd__o221a_1
XPHY_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater651 _14529_/CLK vssd1 vssd1 vccd1 vccd1 _14470_/CLK sky130_fd_sc_hd__buf_8
XFILLER_211_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater662 _14094_/CLK vssd1 vssd1 vccd1 vccd1 _14095_/CLK sky130_fd_sc_hd__buf_12
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _13668_/Q _08792_/X _08556_/X _08793_/X _08794_/X vssd1 vssd1 vccd1 vccd1
+ _13668_/D sky130_fd_sc_hd__o221a_1
XPHY_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater673 _14071_/CLK vssd1 vssd1 vccd1 vccd1 _14119_/CLK sky130_fd_sc_hd__buf_12
Xrepeater684 _12282_/X vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__buf_12
XFILLER_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater695 input39/X vssd1 vssd1 vccd1 vccd1 _12651_/S sky130_fd_sc_hd__buf_4
XPHY_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07747_ _07772_/A vssd1 vssd1 vccd1 vccd1 _07747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07678_ _14223_/Q _07669_/X _07370_/X _07670_/X _07676_/X vssd1 vssd1 vccd1 vccd1
+ _14223_/D sky130_fd_sc_hd__o221a_1
XFILLER_183_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09417_ _09419_/A _13079_/X vssd1 vssd1 vccd1 vccd1 _13320_/D sky130_fd_sc_hd__and2_1
XFILLER_77_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06629_ _06628_/Y _06599_/X _06628_/Y _06599_/X vssd1 vssd1 vccd1 vccd1 _06629_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09348_ _09351_/A _12919_/X vssd1 vssd1 vccd1 vccd1 _13376_/D sky130_fd_sc_hd__and2_1
XFILLER_51_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09279_ _13420_/Q _09275_/X _07708_/A _09277_/X _09267_/X vssd1 vssd1 vccd1 vccd1
+ _13420_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11310_ _11308_/Y _11223_/X _11309_/Y _11225_/X vssd1 vssd1 vccd1 vccd1 _11310_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12290_ _11782_/Y _14553_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__mux2_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ _11239_/Y _11178_/X _11240_/Y _11180_/X vssd1 vssd1 vccd1 vccd1 _11241_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11172_ _11408_/A vssd1 vssd1 vccd1 vccd1 _11172_/X sky130_fd_sc_hd__buf_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _10126_/A _12451_/X vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10054_ _13356_/Q _09970_/B _09971_/A vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__o21a_1
XPHY_7453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13813_ _14123_/CLK _13813_/D vssd1 vssd1 vccd1 vccd1 _13813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13744_ _14130_/CLK _13744_/D vssd1 vssd1 vccd1 vccd1 _13744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10956_ _10939_/Y _10940_/X _10945_/X _10950_/X _10955_/X vssd1 vssd1 vccd1 vccd1
+ _10993_/C sky130_fd_sc_hd__o2111a_4
XFILLER_127_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13675_ _14146_/CLK _13675_/D vssd1 vssd1 vccd1 vccd1 _13675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10887_ _13397_/Q _10804_/X _13709_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _10887_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12626_ _09841_/Y _13331_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__mux2_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12557_ _09954_/X _13302_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11508_ _14080_/Q vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12488_ _12509_/X _06970_/Y _12488_/S vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14227_ _14595_/CLK _14227_/D vssd1 vssd1 vccd1 vccd1 _14227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11439_ _11439_/A vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ _14470_/CLK _14158_/D vssd1 vssd1 vccd1 vccd1 _14158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _12633_/X _13108_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ _14169_/CLK _14089_/D vssd1 vssd1 vccd1 vccd1 _14089_/Q sky130_fd_sc_hd__dfxtp_1
X_06980_ _06974_/X _12315_/X _06979_/Y _06976_/X vssd1 vssd1 vccd1 vccd1 _06981_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08650_ _13747_/Q _08643_/X _08570_/X _08644_/X _08646_/X vssd1 vssd1 vccd1 vccd1
+ _13747_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07601_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07601_/X sky130_fd_sc_hd__clkbuf_2
X_08581_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08581_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07532_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07532_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07463_ _14338_/Q _07459_/X _07377_/X _07460_/X _07461_/X vssd1 vssd1 vccd1 vccd1
+ _14338_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09202_ _09272_/A _11635_/A vssd1 vssd1 vccd1 vccd1 _09258_/A sky130_fd_sc_hd__or2_2
XFILLER_17_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07394_ _08181_/A vssd1 vssd1 vccd1 vccd1 _07394_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09133_ _09189_/A vssd1 vssd1 vccd1 vccd1 _09188_/A sky130_fd_sc_hd__inv_2
XFILLER_13_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09064_ _09132_/A _11660_/A vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__or2_2
XFILLER_198_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08015_ _14056_/Q _07955_/A _07796_/X _07957_/A _08011_/X vssd1 vssd1 vccd1 vccd1
+ _14056_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ _09966_/A vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__inv_2
XFILLER_63_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08917_ _08917_/A vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__buf_6
XFILLER_98_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09897_ _09897_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__or2_1
XPHY_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _13644_/Q _08844_/X _08517_/X _08845_/X _08847_/X vssd1 vssd1 vccd1 vccd1
+ _13644_/D sky130_fd_sc_hd__o221a_1
XFILLER_98_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _13678_/Q _08775_/X _08530_/X _08776_/X _08777_/X vssd1 vssd1 vccd1 vccd1
+ _13678_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10808_/Y _10704_/X _10809_/Y _10706_/X vssd1 vssd1 vccd1 vccd1 _10810_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11790_ _13416_/Q _11747_/X _13735_/Q _12416_/S _11789_/X vssd1 vssd1 vccd1 vccd1
+ _11823_/B sky130_fd_sc_hd__a221oi_2
XPHY_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10741_ _11451_/A vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13460_ _14169_/CLK _13460_/D vssd1 vssd1 vccd1 vccd1 _13460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10672_ _14296_/Q vssd1 vssd1 vccd1 vccd1 _10672_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _13217_/Q _12410_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13391_ _14529_/CLK _13391_/D vssd1 vssd1 vccd1 vccd1 _13391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12342_ _13192_/Q _12341_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12342_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _12063_/Y _13374_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _14130_/CLK _14012_/D vssd1 vssd1 vccd1 vccd1 _14012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11224_ _14463_/Q vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11155_ _14462_/Q vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10106_ _10114_/A _12472_/X vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__nor2_8
XFILLER_1_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11086_ _13954_/Q vssd1 vssd1 vccd1 vccd1 _11086_/Y sky130_fd_sc_hd__inv_2
XPHY_7250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput240 la_oenb[50] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_1
XPHY_7261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 la_oenb[60] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_hd__buf_1
XPHY_7272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10037_ _13374_/Q _10006_/B _10007_/A vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__o21a_1
Xinput262 la_oenb[70] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__buf_1
XFILLER_188_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput273 la_oenb[80] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_hd__buf_1
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput284 la_oenb[90] vssd1 vssd1 vccd1 vccd1 input284/X sky130_fd_sc_hd__buf_1
XPHY_6560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput295 wb_clk_i vssd1 vssd1 vccd1 vccd1 input295/X sky130_fd_sc_hd__buf_4
XFILLER_188_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11988_ _11969_/X _11988_/B _11988_/C _11988_/D vssd1 vssd1 vccd1 vccd1 _11989_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _14047_/CLK _13727_/D vssd1 vssd1 vccd1 vccd1 _13727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ _13951_/Q vssd1 vssd1 vccd1 vccd1 _10939_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13658_ _14047_/CLK _13658_/D vssd1 vssd1 vccd1 vccd1 _13658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _09854_/Y _13324_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12609_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13589_ _14183_/CLK _13589_/D vssd1 vssd1 vccd1 vccd1 _13589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _09820_/A vssd1 vssd1 vccd1 vccd1 _09820_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09751_ _13337_/Q vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__inv_2
XFILLER_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06963_ _06972_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _14572_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08702_ _13721_/Q _08698_/X _08519_/X _08699_/X _08696_/X vssd1 vssd1 vccd1 vccd1
+ _13721_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09682_ _06869_/A _09610_/A _14596_/Q _09610_/Y vssd1 vssd1 vccd1 vccd1 _09682_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06894_ _06880_/X _12292_/X _06893_/X _06883_/X vssd1 vssd1 vccd1 vccd1 _06895_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_67_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _13756_/Q _08626_/X _08632_/X _08627_/X _08628_/X vssd1 vssd1 vccd1 vccd1
+ _13756_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _13789_/Q _08552_/X _08562_/X _08554_/X _08563_/X vssd1 vssd1 vccd1 vccd1
+ _13789_/D sky130_fd_sc_hd__o221a_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07515_ _14311_/Q _07508_/X _07345_/X _07509_/X _07511_/X vssd1 vssd1 vccd1 vccd1
+ _14311_/D sky130_fd_sc_hd__o221a_1
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08495_ _13815_/Q _08486_/X _08494_/X _08488_/X _08480_/X vssd1 vssd1 vccd1 vccd1
+ _13815_/D sky130_fd_sc_hd__o221a_1
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07446_ _14348_/Q _07440_/X _07352_/X _07441_/X _07444_/X vssd1 vssd1 vccd1 vccd1
+ _14348_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07377_ _08165_/A vssd1 vssd1 vccd1 vccd1 _07377_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09116_ _13510_/Q _09111_/X _08965_/X _09112_/X _09109_/X vssd1 vssd1 vccd1 vccd1
+ _13510_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09047_ _13548_/Q _09039_/X _08967_/X _09040_/X _09045_/X vssd1 vssd1 vccd1 vccd1
+ _13548_/D sky130_fd_sc_hd__o221a_1
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12960_ _12560_/X input335/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _13653_/Q vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__inv_2
XPHY_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12533_/X _12890_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14633_/CLK _14630_/D vssd1 vssd1 vccd1 vccd1 _14630_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11842_ _13534_/Q vssd1 vssd1 vccd1 vccd1 _11842_/Y sky130_fd_sc_hd__inv_2
XPHY_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14595_/CLK _14561_/D vssd1 vssd1 vccd1 vccd1 _14561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11773_ _11771_/Y _11683_/X _11772_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11773_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _14110_/CLK _13512_/D vssd1 vssd1 vccd1 vccd1 _13512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _14492_/Q vssd1 vssd1 vccd1 vccd1 _10724_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14495_/CLK _14492_/D vssd1 vssd1 vccd1 vccd1 _14492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13443_ _14459_/CLK _13443_/D vssd1 vssd1 vccd1 vccd1 _13443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10655_ _13867_/Q vssd1 vssd1 vccd1 vccd1 _10655_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13374_ _14573_/CLK _13374_/D vssd1 vssd1 vccd1 vccd1 _13374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10586_ _14606_/Q vssd1 vssd1 vccd1 vccd1 _10586_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ _12324_/X _13198_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12325_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12256_ _12040_/Y _13357_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12256_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11207_ _11198_/Y _11199_/X _11200_/Y _11201_/X _11206_/X vssd1 vssd1 vccd1 vccd1
+ _11228_/B sky130_fd_sc_hd__o221a_1
XFILLER_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ vssd1 vssd1 vccd1 vccd1 _12187_/HI _12187_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11138_ _13558_/Q _10958_/X _13799_/Q _10959_/X vssd1 vssd1 vccd1 vccd1 _11138_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11069_ _11064_/Y _10973_/X _11065_/Y _10975_/X _11068_/X vssd1 vssd1 vccd1 vccd1
+ _11076_/C sky130_fd_sc_hd__o221a_1
XPHY_7080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07300_ _14405_/Q _07238_/A _06850_/B _07240_/A _07295_/X vssd1 vssd1 vccd1 vccd1
+ _14405_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08280_ _13933_/Q _08274_/X _08101_/X _08276_/X _08278_/X vssd1 vssd1 vccd1 vccd1
+ _13933_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07231_ _09272_/A vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__buf_2
XFILLER_144_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07162_ _07218_/A vssd1 vssd1 vccd1 vccd1 _07217_/A sky130_fd_sc_hd__inv_2
XFILLER_146_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07093_ _07145_/A vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput500 _12131_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__clkbuf_2
Xoutput511 _12141_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput522 _12151_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput533 _12161_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput544 _12171_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__clkbuf_2
Xoutput555 _12181_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__clkbuf_2
Xoutput566 _12191_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput577 _13265_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput588 _13275_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput599 _13285_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_2
X_09803_ _09801_/A _09801_/B _09802_/Y vssd1 vssd1 vccd1 vccd1 _09803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _08017_/A vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _12603_/S vssd1 vssd1 vccd1 vccd1 _12232_/A sky130_fd_sc_hd__clkinv_16
XFILLER_189_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06946_ _14576_/Q vssd1 vssd1 vccd1 vccd1 _06946_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _12667_/S vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__inv_2
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06877_ _06877_/A _06877_/B vssd1 vssd1 vccd1 vccd1 _14594_/D sky130_fd_sc_hd__nor2_1
X_08616_ _13766_/Q _08610_/X _08521_/X _08611_/X _08612_/X vssd1 vssd1 vccd1 vccd1
+ _13766_/D sky130_fd_sc_hd__o221a_1
XFILLER_76_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09596_ _09557_/A _09595_/X _13256_/Q _09545_/A vssd1 vssd1 vccd1 vccd1 _13224_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _13796_/Q _08540_/X _08546_/X _08542_/X _08538_/X vssd1 vssd1 vccd1 vccd1
+ _13796_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08478_ _13821_/Q _08415_/A _08188_/X _08417_/A _08474_/X vssd1 vssd1 vccd1 vccd1
+ _13821_/D sky130_fd_sc_hd__o221a_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07429_ _14357_/Q _07422_/X _07428_/X _07424_/X _07425_/X vssd1 vssd1 vccd1 vccd1
+ _14357_/D sky130_fd_sc_hd__o221a_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10440_ _11408_/A vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _14251_/Q vssd1 vssd1 vccd1 vccd1 _10371_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ vssd1 vssd1 vccd1 vccd1 _12110_/HI _12110_/LO sky130_fd_sc_hd__conb_1
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13090_ _13089_/X _12623_/X _13110_/S vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12041_ _09776_/A _12035_/X _09888_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12041_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_65_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13992_ _14107_/CLK _13992_/D vssd1 vssd1 vccd1 vccd1 _13992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12943_ _12551_/X _12942_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_120 _10838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _12529_/X _12873_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11825_ _13456_/Q vssd1 vssd1 vccd1 vccd1 _11825_/Y sky130_fd_sc_hd__inv_2
XANTENNA_153 _11865_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14627_/CLK _14613_/D vssd1 vssd1 vccd1 vccd1 _14613_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_164 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 input332/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 input344/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 input358/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544_ _14621_/CLK _14544_/D vssd1 vssd1 vccd1 vccd1 _14544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11756_ _11754_/Y _11653_/X _11755_/Y _11655_/X vssd1 vssd1 vccd1 vccd1 _11756_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ _10703_/Y _10704_/X _10705_/Y _10706_/X vssd1 vssd1 vccd1 vccd1 _10707_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14475_ _14527_/CLK _14475_/D vssd1 vssd1 vccd1 vccd1 _14475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11678_/Y _11679_/X _11680_/Y _11681_/X _11686_/X vssd1 vssd1 vccd1 vccd1
+ _11698_/C sky130_fd_sc_hd__o221a_1
XFILLER_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13426_ _14139_/CLK _13426_/D vssd1 vssd1 vccd1 vccd1 _13426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10638_ _14139_/Q vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13357_ _14639_/CLK _13357_/D vssd1 vssd1 vccd1 vccd1 _13357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10569_ _13390_/Q _10568_/X _13702_/Q _10440_/X vssd1 vssd1 vccd1 vccd1 _10569_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12308_ _10921_/Y _14535_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13288_ _13996_/CLK _13288_/D vssd1 vssd1 vccd1 vccd1 _13288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12239_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06800_ _08954_/A vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__buf_2
XFILLER_81_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07780_ _08171_/A vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__buf_4
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XFILLER_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06731_ _14633_/Q _06530_/X _06725_/X _06726_/X _06730_/X vssd1 vssd1 vccd1 vccd1
+ _14633_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09450_ _09450_/A _12931_/X vssd1 vssd1 vccd1 vccd1 _13293_/D sky130_fd_sc_hd__and2_1
X_06662_ _06655_/X _06661_/Y _06655_/X _06661_/Y vssd1 vssd1 vccd1 vccd1 _06662_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08401_ _13864_/Q _08396_/X _08179_/X _08397_/X _08400_/X vssd1 vssd1 vccd1 vccd1
+ _13864_/D sky130_fd_sc_hd__o221a_1
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09381_ _09382_/A _13155_/X vssd1 vssd1 vccd1 vccd1 _13349_/D sky130_fd_sc_hd__and2_1
XFILLER_55_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06593_ _06595_/A vssd1 vssd1 vccd1 vccd1 _06593_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08332_ _13902_/Q _08326_/X _08181_/X _08327_/X _08329_/X vssd1 vssd1 vccd1 vccd1
+ _13902_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08263_ _13940_/Q _08255_/X _08183_/X _08256_/X _08257_/X vssd1 vssd1 vccd1 vccd1
+ _13940_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07214_ _14454_/Q _07209_/X _06814_/X _07210_/X _07213_/X vssd1 vssd1 vccd1 vccd1
+ _14454_/D sky130_fd_sc_hd__o221a_1
X_08194_ _08814_/A _08340_/B _08814_/C _08584_/D vssd1 vssd1 vccd1 vccd1 _11646_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ _07145_/A vssd1 vssd1 vccd1 vccd1 _07145_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07076_ _14526_/Q _07069_/X _06834_/X _07070_/X _07071_/X vssd1 vssd1 vccd1 vccd1
+ _14526_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput374 _12211_/X vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput385 _12221_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput396 _12231_/X vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07978_/X sky130_fd_sc_hd__buf_2
XFILLER_19_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ _09715_/X _09716_/X _09715_/X _09716_/X vssd1 vssd1 vccd1 vccd1 _09717_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06929_ _06935_/A _06929_/B vssd1 vssd1 vccd1 vccd1 _14581_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _09628_/X _09647_/Y _09628_/X _09647_/Y vssd1 vssd1 vccd1 vccd1 _09648_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09570_/X _09578_/X _13263_/Q _09571_/X vssd1 vssd1 vccd1 vccd1 _13231_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _13568_/Q _11430_/X _13809_/Q _11431_/X vssd1 vssd1 vccd1 vccd1 _11610_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _13318_/Q _12589_/X _12655_/S vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__mux2_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11536_/Y _11445_/X _11537_/Y _11447_/X _11540_/X vssd1 vssd1 vccd1 vccd1
+ _11548_/C sky130_fd_sc_hd__o221a_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _14305_/CLK _14260_/D vssd1 vssd1 vccd1 vccd1 _14260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11472_ _13409_/Q _11278_/X _13721_/Q _11408_/X vssd1 vssd1 vccd1 vccd1 _11472_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ _13368_/CLK _13211_/D vssd1 vssd1 vccd1 vccd1 _13211_/Q sky130_fd_sc_hd__dfxtp_2
X_10423_ _14058_/Q vssd1 vssd1 vccd1 vccd1 _10423_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14191_ _14305_/CLK _14191_/D vssd1 vssd1 vccd1 vccd1 _14191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13142_ _13141_/X _12649_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _14095_/Q vssd1 vssd1 vccd1 vccd1 _10354_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13073_ _12616_/X _13072_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__mux2_1
X_10285_ _14288_/Q vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12024_ _14169_/Q vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13975_ _14095_/CLK _13975_/D vssd1 vssd1 vccd1 vccd1 _13975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ _12925_/X _12543_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _12525_/X _12856_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11808_ _11806_/Y _11673_/X _11807_/Y _11675_/X vssd1 vssd1 vccd1 vccd1 _11808_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12788_ _09533_/X input347/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11739_ _11720_/X _11739_/B _11739_/C _11739_/D vssd1 vssd1 vccd1 vccd1 _11740_/D
+ sky130_fd_sc_hd__and4b_1
X_14527_ _14527_/CLK _14527_/D vssd1 vssd1 vccd1 vccd1 _14527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14458_ _14595_/CLK _14458_/D vssd1 vssd1 vccd1 vccd1 _14458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13409_ _14183_/CLK _13409_/D vssd1 vssd1 vccd1 vccd1 _13409_/Q sky130_fd_sc_hd__dfxtp_1
X_14389_ _14629_/CLK _14389_/D vssd1 vssd1 vccd1 vccd1 _14389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08950_ _08950_/A vssd1 vssd1 vccd1 vccd1 _08950_/X sky130_fd_sc_hd__buf_4
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07901_ _14121_/Q _07892_/X _07728_/X _07894_/X _07897_/X vssd1 vssd1 vccd1 vccd1
+ _14121_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08881_ _13624_/Q _08876_/X _08648_/X _08877_/X _08880_/X vssd1 vssd1 vccd1 vccd1
+ _13624_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07832_ _14159_/Q _07829_/X _07733_/X _07830_/X _07831_/X vssd1 vssd1 vccd1 vccd1
+ _14159_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07763_ _14187_/Q _07758_/X _07762_/X _07760_/X _07756_/X vssd1 vssd1 vccd1 vccd1
+ _14187_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09502_ _13261_/Q _09500_/X _12256_/X _09501_/X vssd1 vssd1 vccd1 vccd1 _13261_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06714_ _07708_/A vssd1 vssd1 vccd1 vccd1 _06714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07694_ _14213_/Q _07687_/X _07396_/X _07688_/X _07692_/X vssd1 vssd1 vccd1 vccd1
+ _14213_/D sky130_fd_sc_hd__o221a_1
XFILLER_183_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09433_ _09445_/A vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__buf_2
XFILLER_77_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06645_ _06668_/A vssd1 vssd1 vccd1 vccd1 _06645_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09364_ _09364_/A _12843_/X vssd1 vssd1 vccd1 vccd1 _13363_/D sky130_fd_sc_hd__and2_1
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06576_ input94/X vssd1 vssd1 vccd1 vccd1 _08977_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08315_ _13913_/Q _08310_/X _08155_/X _08311_/X _08313_/X vssd1 vssd1 vccd1 vccd1
+ _13913_/D sky130_fd_sc_hd__o221a_1
XFILLER_205_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_20 _11989_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_31 _08243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _07367_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08246_ _08246_/A vssd1 vssd1 vccd1 vccd1 _08246_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_53 _07764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 _07872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_75 _08171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_86 _08606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_97 _08967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08177_ _13983_/Q _08174_/X _08175_/X _08176_/X _08172_/X vssd1 vssd1 vccd1 vccd1
+ _13983_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07128_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07059_ _14536_/Q _07052_/X _07058_/X _07053_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _14536_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10070_ _10070_/A _12507_/S vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__or2_2
XFILLER_173_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13760_ _13996_/CLK _13760_/D vssd1 vssd1 vccd1 vccd1 _13760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10972_ _14302_/Q vssd1 vssd1 vccd1 vccd1 _10972_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12711_ _09565_/X _12710_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13204_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13691_ _14056_/CLK _13691_/D vssd1 vssd1 vccd1 vccd1 _13691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12642_ _09828_/Y _13339_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12642_/X sky130_fd_sc_hd__mux2_1
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _09942_/X _13310_/Q _12603_/S vssd1 vssd1 vccd1 vccd1 _12573_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ _14527_/CLK _14312_/D vssd1 vssd1 vccd1 vccd1 _14312_/Q sky130_fd_sc_hd__dfxtp_1
X_11524_ _14002_/Q vssd1 vssd1 vccd1 vccd1 _11524_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _14325_/CLK _14243_/D vssd1 vssd1 vccd1 vccd1 _14243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11455_ _11455_/A vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ _14369_/Q vssd1 vssd1 vccd1 vccd1 _10406_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14174_ _14178_/CLK _14174_/D vssd1 vssd1 vccd1 vccd1 _14174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _11384_/Y _11213_/X _11385_/Y _11215_/X vssd1 vssd1 vccd1 vccd1 _11386_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13125_ _12641_/X _13124_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__mux2_1
X_10337_ _10335_/Y _10248_/X _10336_/Y _10251_/X vssd1 vssd1 vccd1 vccd1 _10337_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13056_ _12608_/X input358/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__mux2_1
X_10268_ _13820_/Q vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12007_ _12005_/Y _10195_/A _12006_/Y _10198_/A vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _10193_/Y _10195_/X _10196_/Y _10198_/X vssd1 vssd1 vccd1 vccd1 _10199_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13958_ _13996_/CLK _13958_/D vssd1 vssd1 vccd1 vccd1 _13958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12909_ _12538_/X _12908_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ _14100_/CLK _13889_/D vssd1 vssd1 vccd1 vccd1 _13889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08100_ _14012_/Q _08095_/X _08099_/X _08097_/X _08089_/X vssd1 vssd1 vccd1 vccd1
+ _14012_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09080_ _13533_/Q _09077_/X _08833_/X _09079_/X _09074_/X vssd1 vssd1 vccd1 vccd1
+ _13533_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08031_ _08133_/A vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__buf_2
Xinput40 la_data_in[100] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
XFILLER_15_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 la_data_in[110] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_1
XFILLER_190_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput62 la_data_in[120] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_1
XFILLER_176_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput73 la_data_in[15] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_1
Xinput84 la_data_in[25] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_1
XFILLER_196_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput95 la_data_in[35] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09982_ _13362_/Q _09982_/B vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08933_ _08933_/A vssd1 vssd1 vccd1 vccd1 _08933_/X sky130_fd_sc_hd__buf_6
XFILLER_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08864_ _13634_/Q _08860_/X _08544_/X _08861_/X _08863_/X vssd1 vssd1 vccd1 vccd1
+ _13634_/D sky130_fd_sc_hd__o221a_1
XPHY_6219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater630 _10097_/A vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07815_ _14167_/Q _07808_/X _07710_/X _07811_/X _07812_/X vssd1 vssd1 vccd1 vccd1
+ _14167_/D sky130_fd_sc_hd__o221a_1
XPHY_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater641 _14459_/CLK vssd1 vssd1 vccd1 vccd1 _14595_/CLK sky130_fd_sc_hd__buf_12
Xrepeater652 _14481_/CLK vssd1 vssd1 vccd1 vccd1 _14325_/CLK sky130_fd_sc_hd__buf_12
X_08795_ _13669_/Q _08792_/X _08553_/X _08793_/X _08794_/X vssd1 vssd1 vccd1 vccd1
+ _13669_/D sky130_fd_sc_hd__o221a_1
Xrepeater663 _14123_/CLK vssd1 vssd1 vccd1 vccd1 _14130_/CLK sky130_fd_sc_hd__buf_12
XPHY_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater674 _13877_/CLK vssd1 vssd1 vccd1 vccd1 _14639_/CLK sky130_fd_sc_hd__buf_12
XFILLER_42_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater685 _12396_/S vssd1 vssd1 vccd1 vccd1 _12417_/S sky130_fd_sc_hd__buf_8
XPHY_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07746_ _08137_/A vssd1 vssd1 vccd1 vccd1 _07746_/X sky130_fd_sc_hd__buf_6
XPHY_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater696 _13121_/S vssd1 vssd1 vccd1 vccd1 _13177_/S sky130_fd_sc_hd__buf_8
XFILLER_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07677_ _14224_/Q _07669_/X _07456_/X _07670_/X _07676_/X vssd1 vssd1 vccd1 vccd1
+ _14224_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09416_ _09419_/A _13075_/X vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__and2_1
XFILLER_73_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06628_ input99/X vssd1 vssd1 vccd1 vccd1 _06628_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09347_ _09351_/A _12915_/X vssd1 vssd1 vccd1 vccd1 _13377_/D sky130_fd_sc_hd__and2_1
XFILLER_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06559_ _06559_/A vssd1 vssd1 vccd1 vccd1 _06559_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09278_ _13421_/Q _09275_/X _07809_/A _09277_/X _09267_/X vssd1 vssd1 vccd1 vccd1
+ _13421_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08229_ _08246_/A vssd1 vssd1 vccd1 vccd1 _08229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11240_ _13879_/Q vssd1 vssd1 vccd1 vccd1 _11240_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11171_ _11407_/A vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_190_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10122_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _12449_/S sky130_fd_sc_hd__or2_1
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10053_ _13355_/Q _10052_/A _09969_/A vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__o21a_1
XPHY_7443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13812_ _14123_/CLK _13812_/D vssd1 vssd1 vccd1 vccd1 _13812_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13743_ _14130_/CLK _13743_/D vssd1 vssd1 vccd1 vccd1 _13743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10955_ _10951_/Y _10952_/X _10953_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _10955_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13674_ _14071_/CLK _13674_/D vssd1 vssd1 vccd1 vccd1 _13674_/Q sky130_fd_sc_hd__dfxtp_1
X_10886_ _10881_/Y _10687_/X _10882_/Y _10689_/X _10885_/X vssd1 vssd1 vccd1 vccd1
+ _10921_/A sky130_fd_sc_hd__o221a_2
XFILLER_38_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12625_ _13332_/Q _12624_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__mux2_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ _13287_/Q _09955_/X _12619_/S vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11507_ _11507_/A _11507_/B _11507_/C _11507_/D vssd1 vssd1 vccd1 vccd1 _11507_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12486_/X _06967_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12487_/X sky130_fd_sc_hd__mux2_2
XFILLER_176_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11438_ _14624_/Q vssd1 vssd1 vccd1 vccd1 _11438_/Y sky130_fd_sc_hd__inv_2
X_14226_ _14459_/CLK _14226_/D vssd1 vssd1 vccd1 vccd1 _14226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _14305_/CLK _14157_/D vssd1 vssd1 vccd1 vccd1 _14157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11369_ _11367_/Y _11183_/X _11368_/Y _11185_/X vssd1 vssd1 vccd1 vccd1 _11369_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ _12633_/X input361/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14088_ _14169_/CLK _14088_/D vssd1 vssd1 vccd1 vccd1 _14088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13039_ _12598_/X _13038_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07600_ _14265_/Q _07597_/X _07365_/X _07598_/X _07593_/X vssd1 vssd1 vccd1 vccd1
+ _14265_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08580_ _13782_/Q _08486_/A _08579_/X _08488_/A _08575_/X vssd1 vssd1 vccd1 vccd1
+ _13782_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ _14301_/Q _07524_/X _07370_/X _07525_/X _07527_/X vssd1 vssd1 vccd1 vccd1
+ _14301_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07462_ _14339_/Q _07459_/X _07374_/X _07460_/X _07461_/X vssd1 vssd1 vccd1 vccd1
+ _14339_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09201_ _09271_/A _09201_/B _09201_/C _09201_/D vssd1 vssd1 vccd1 vccd1 _11635_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07393_ _14371_/Q _07387_/X _07392_/X _07389_/X _07385_/X vssd1 vssd1 vccd1 vccd1
+ _14371_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09132_ _09132_/A _11693_/A vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__or2_2
XFILLER_194_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _09271_/A _09063_/B _09063_/C _09201_/D vssd1 vssd1 vccd1 vccd1 _11660_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_15_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08014_ _14057_/Q _08007_/X _07792_/X _08008_/X _08011_/X vssd1 vssd1 vccd1 vccd1
+ _14057_/D sky130_fd_sc_hd__o221a_1
XFILLER_102_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09965_ _13352_/Q _13351_/Q vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__nand2_4
XFILLER_115_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08916_ _08956_/A vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _09896_/A _09952_/A vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__or2_2
XFILLER_44_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08871_/A vssd1 vssd1 vccd1 vccd1 _08847_/X sky130_fd_sc_hd__buf_2
XPHY_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ _13679_/Q _08775_/X _08527_/X _08776_/X _08777_/X vssd1 vssd1 vccd1 vccd1
+ _13679_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__buf_2
XPHY_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _14258_/Q vssd1 vssd1 vccd1 vccd1 _10740_/Y sky130_fd_sc_hd__inv_2
XPHY_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10671_ _10666_/Y _10478_/X _10667_/Y _10481_/X _10670_/X vssd1 vssd1 vccd1 vccd1
+ _10684_/B sky130_fd_sc_hd__o221a_4
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _13217_/Q _06696_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12410_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13390_ _14529_/CLK _13390_/D vssd1 vssd1 vccd1 vccd1 _13390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12341_ _13192_/Q _06850_/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ _12062_/Y _13373_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12272_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14011_ _14130_/CLK _14011_/D vssd1 vssd1 vccd1 vccd1 _14011_/Q sky130_fd_sc_hd__dfxtp_1
X_11223_ _11459_/A vssd1 vssd1 vccd1 vccd1 _11223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11154_ _13480_/Q vssd1 vssd1 vccd1 vccd1 _11154_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10105_ _10141_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _12470_/S sky130_fd_sc_hd__or2_1
XFILLER_150_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11085_ _14227_/Q _10933_/X _14422_/Q _10935_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11118_/B sky130_fd_sc_hd__a221oi_2
XPHY_7240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput230 la_oenb[41] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_1
XFILLER_62_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput241 la_oenb[51] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_1
XFILLER_23_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ _13373_/Q _10004_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _10036_/X sky130_fd_sc_hd__o21a_1
Xinput252 la_oenb[61] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__buf_1
XFILLER_0_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput263 la_oenb[71] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_hd__buf_1
XPHY_7284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput274 la_oenb[81] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_hd__buf_1
XPHY_7295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput285 la_oenb[91] vssd1 vssd1 vccd1 vccd1 input285/X sky130_fd_sc_hd__buf_1
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput296 wb_rst_i vssd1 vssd1 vccd1 vccd1 input296/X sky130_fd_sc_hd__buf_4
XPHY_6572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11987_ _11982_/Y _10242_/A _11983_/Y _10245_/A _11986_/X vssd1 vssd1 vccd1 vccd1
+ _11988_/D sky130_fd_sc_hd__o221a_1
XPHY_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13726_ _14178_/CLK _13726_/D vssd1 vssd1 vccd1 vccd1 _13726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10938_ _14224_/Q _10933_/X _14419_/Q _10935_/X _10937_/X vssd1 vssd1 vccd1 vccd1
+ _10993_/B sky130_fd_sc_hd__a221oi_2
XFILLER_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13657_ _14056_/CLK _13657_/D vssd1 vssd1 vccd1 vccd1 _13657_/Q sky130_fd_sc_hd__dfxtp_1
X_10869_ _14183_/Q vssd1 vssd1 vccd1 vccd1 _10869_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _13325_/Q _12607_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _14188_/CLK _13588_/D vssd1 vssd1 vccd1 vccd1 _13588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ _13377_/Q _10015_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12539_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14209_ _14325_/CLK _14209_/D vssd1 vssd1 vccd1 vccd1 _14209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _13338_/Q vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__inv_2
X_06962_ _06956_/X _12310_/X _06961_/Y _06958_/X vssd1 vssd1 vccd1 vccd1 _06963_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08701_ _13722_/Q _08698_/X _08517_/X _08699_/X _08696_/X vssd1 vssd1 vccd1 vccd1
+ _13722_/D sky130_fd_sc_hd__o221a_1
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _12507_/S sky130_fd_sc_hd__buf_6
XFILLER_132_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06893_ _06893_/A vssd1 vssd1 vccd1 vccd1 _06893_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08632_ _09035_/A vssd1 vssd1 vccd1 vccd1 _08632_/X sky130_fd_sc_hd__buf_4
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08563_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08563_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07514_ _14312_/Q _07508_/X _07343_/X _07509_/X _07511_/X vssd1 vssd1 vccd1 vccd1
+ _14312_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08494_ _08827_/A vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07445_ _14349_/Q _07440_/X _07349_/X _07441_/X _07444_/X vssd1 vssd1 vccd1 vccd1
+ _14349_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07376_ _14378_/Q _07373_/X _07374_/X _07375_/X _07371_/X vssd1 vssd1 vccd1 vccd1
+ _14378_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09115_ _13511_/Q _09111_/X _08962_/X _09112_/X _09109_/X vssd1 vssd1 vccd1 vccd1
+ _13511_/D sky130_fd_sc_hd__o221a_1
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _13549_/Q _09039_/X _08965_/X _09040_/X _09045_/X vssd1 vssd1 vccd1 vccd1
+ _13549_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09948_ _13298_/Q _09946_/Y _09893_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09879_ _13289_/Q vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__inv_2
XFILLER_115_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11910_ _13692_/Q vssd1 vssd1 vccd1 vccd1 _11910_/Y sky130_fd_sc_hd__inv_2
XPHY_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12533_/X _12889_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12890_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11841_ _14009_/Q vssd1 vssd1 vccd1 vccd1 _11841_/Y sky130_fd_sc_hd__inv_2
XPHY_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11772_ _14280_/Q vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__inv_2
XPHY_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14595_/CLK _14560_/D vssd1 vssd1 vccd1 vccd1 _14560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _13201_/Q _10539_/X _14024_/Q _10719_/X _10722_/X vssd1 vssd1 vccd1 vccd1
+ _10723_/X sky130_fd_sc_hd__a221o_2
X_13511_ _14110_/CLK _13511_/D vssd1 vssd1 vccd1 vccd1 _13511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _14495_/CLK _14491_/D vssd1 vssd1 vccd1 vccd1 _14491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10654_ _13750_/Q vssd1 vssd1 vccd1 vccd1 _10654_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13442_ _14459_/CLK _13442_/D vssd1 vssd1 vccd1 vccd1 _13442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13373_ _14573_/CLK _13373_/D vssd1 vssd1 vccd1 vccd1 _13373_/Q sky130_fd_sc_hd__dfxtp_1
X_10585_ _14333_/Q vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ _13198_/Q _12323_/X input78/X vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12255_ _12039_/Y _13356_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12255_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11206_ _11202_/Y _11203_/X _11204_/Y _11205_/X vssd1 vssd1 vccd1 vccd1 _11206_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12186_ vssd1 vssd1 vccd1 vccd1 _12186_/HI _12186_/LO sky130_fd_sc_hd__conb_1
XFILLER_116_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11137_ _11127_/Y _10940_/X _11130_/X _11133_/X _11136_/X vssd1 vssd1 vccd1 vccd1
+ _11159_/C sky130_fd_sc_hd__o2111a_4
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11068_ _11066_/Y _10977_/X _11067_/Y _10979_/X vssd1 vssd1 vccd1 vccd1 _11068_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _10019_/A vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__inv_2
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13709_ _14146_/CLK _13709_/D vssd1 vssd1 vccd1 vccd1 _13709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _14443_/Q _07164_/A _07083_/X _07166_/A _07228_/X vssd1 vssd1 vccd1 vccd1
+ _14443_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07161_ _08660_/A _11695_/A vssd1 vssd1 vccd1 vccd1 _07218_/A sky130_fd_sc_hd__or2_2
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07092_ _07092_/A vssd1 vssd1 vccd1 vccd1 _07092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput501 _12132_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput512 _12142_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__clkbuf_2
Xoutput523 _12152_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput534 _12162_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__clkbuf_2
Xoutput545 _12172_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput556 _12182_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__clkbuf_2
Xoutput567 _12192_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput578 _13266_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput589 _13276_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09802_ _09805_/B vssd1 vssd1 vccd1 vccd1 _09802_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07994_ _14070_/Q _07991_/X _07762_/X _07992_/X _07987_/X vssd1 vssd1 vccd1 vccd1
+ _14070_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09733_ _09733_/A vssd1 vssd1 vccd1 vccd1 _12509_/S sky130_fd_sc_hd__clkbuf_2
X_06945_ _06954_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _14577_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09664_ _10060_/A vssd1 vssd1 vccd1 vccd1 _12506_/S sky130_fd_sc_hd__clkinv_8
X_06876_ _06857_/X _12288_/X _06875_/Y _06861_/X vssd1 vssd1 vccd1 vccd1 _06877_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _13767_/Q _08610_/X _08519_/X _08611_/X _08612_/X vssd1 vssd1 vccd1 vccd1
+ _13767_/D sky130_fd_sc_hd__o221a_1
X_09595_ _09597_/A _12343_/X vssd1 vssd1 vccd1 vccd1 _09595_/X sky130_fd_sc_hd__and2_1
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08950_/A vssd1 vssd1 vccd1 vccd1 _08546_/X sky130_fd_sc_hd__buf_4
XFILLER_70_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08477_ _13822_/Q _08415_/A _08186_/X _08417_/A _08474_/X vssd1 vssd1 vccd1 vccd1
+ _13822_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ _08217_/A vssd1 vssd1 vccd1 vccd1 _07428_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07359_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10370_ _14173_/Q vssd1 vssd1 vccd1 vccd1 _10370_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09029_ _13558_/Q _09022_/X _08942_/X _09023_/X _09027_/X vssd1 vssd1 vccd1 vccd1
+ _13558_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _09775_/A _12035_/X _09887_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12040_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _14107_/CLK _13991_/D vssd1 vssd1 vccd1 vccd1 _13991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12942_ _12941_/X _12551_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_110 _11449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ _12529_/X _12872_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12873_/X sky130_fd_sc_hd__mux2_1
XPHY_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _10838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_132 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14612_ _14627_/CLK _14612_/D vssd1 vssd1 vccd1 vccd1 _14612_/Q sky130_fd_sc_hd__dfxtp_1
X_11824_ _14087_/Q vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__inv_2
XPHY_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_154 _11887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_165 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 input332/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_187 input348/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 input361/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ _14621_/CLK _14543_/D vssd1 vssd1 vccd1 vccd1 _14543_/Q sky130_fd_sc_hd__dfxtp_1
X_11755_ _14124_/Q vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _11416_/A vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14474_ _14527_/CLK _14474_/D vssd1 vssd1 vccd1 vccd1 _14474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11686_ _11682_/Y _11683_/X _11684_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11686_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ _14056_/CLK _13425_/D vssd1 vssd1 vccd1 vccd1 _13425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10637_ _13905_/Q vssd1 vssd1 vccd1 vccd1 _10637_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10568_ _11042_/A vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__clkbuf_2
X_13356_ _14639_/CLK _13356_/D vssd1 vssd1 vccd1 vccd1 _13356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _10993_/Y _14536_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12307_/X sky130_fd_sc_hd__mux2_2
XFILLER_143_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10499_ _14253_/Q vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__inv_2
X_13287_ _13996_/CLK _13287_/D vssd1 vssd1 vccd1 vccd1 _13287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12238_ _12238_/A vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ vssd1 vssd1 vccd1 vccd1 _12169_/HI _12169_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_06730_ _06785_/A vssd1 vssd1 vccd1 vccd1 _06730_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06661_ _06658_/X _06660_/X _06658_/X _06660_/X vssd1 vssd1 vccd1 vccd1 _06661_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_149_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08400_ _08421_/A vssd1 vssd1 vccd1 vccd1 _08400_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09380_ _09382_/A _13151_/X vssd1 vssd1 vccd1 vccd1 _13350_/D sky130_fd_sc_hd__and2_1
XFILLER_94_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06592_ _06588_/Y _06589_/Y _08967_/A _08974_/A vssd1 vssd1 vccd1 vccd1 _06592_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ _13903_/Q _08326_/X _08179_/X _08327_/X _08329_/X vssd1 vssd1 vccd1 vccd1
+ _13903_/D sky130_fd_sc_hd__o221a_1
XFILLER_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08262_ _13941_/Q _08255_/X _08181_/X _08256_/X _08257_/X vssd1 vssd1 vccd1 vccd1
+ _13941_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07213_ _07213_/A vssd1 vssd1 vccd1 vccd1 _07213_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08193_ _08482_/D vssd1 vssd1 vccd1 vccd1 _08584_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_140_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07144_ _07144_/A vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07075_ _14527_/Q _07069_/X _06831_/X _07070_/X _07071_/X vssd1 vssd1 vccd1 vccd1
+ _14527_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput375 _12212_/X vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput386 _12222_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput397 _12231_/A vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07977_ _14080_/Q _07974_/X _07736_/X _07975_/X _07970_/X vssd1 vssd1 vccd1 vccd1
+ _14080_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09716_ _06924_/Y _06930_/Y _14582_/Q _14580_/Q vssd1 vssd1 vccd1 vccd1 _09716_/X
+ sky130_fd_sc_hd__a22o_1
X_06928_ _06919_/X _12301_/X _06927_/Y _06921_/X vssd1 vssd1 vccd1 vccd1 _06929_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09647_ _09635_/X _09646_/X _09635_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _09647_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06859_ _12417_/S _09650_/A vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__or2_1
XFILLER_3_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ _09586_/A _12370_/X vssd1 vssd1 vccd1 vccd1 _09578_/X sky130_fd_sc_hd__and2_1
XFILLER_73_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _13803_/Q _08526_/X _08527_/X _08528_/X _08524_/X vssd1 vssd1 vccd1 vccd1
+ _13803_/D sky130_fd_sc_hd__o221a_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11540_ _11538_/Y _11449_/X _11539_/Y _11451_/X vssd1 vssd1 vccd1 vccd1 _11540_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11471_ _11466_/Y _11397_/X _11467_/Y _11399_/X _11470_/X vssd1 vssd1 vccd1 vccd1
+ _11507_/A sky130_fd_sc_hd__o221a_2
XFILLER_13_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10422_ _10422_/A _10422_/B _10422_/C _10422_/D vssd1 vssd1 vccd1 vccd1 _10422_/Y
+ sky130_fd_sc_hd__nand4_4
X_13210_ _13368_/CLK _13210_/D vssd1 vssd1 vccd1 vccd1 _13210_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14190_ _14305_/CLK _14190_/D vssd1 vssd1 vccd1 vccd1 _14190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10353_ _13822_/Q vssd1 vssd1 vccd1 vccd1 _10353_/Y sky130_fd_sc_hd__inv_2
X_13141_ _12649_/X _13140_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13072_ _12616_/X input352/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__mux2_1
X_10284_ _10279_/Y _10214_/X _10280_/Y _10217_/X _10283_/X vssd1 vssd1 vccd1 vccd1
+ _10297_/B sky130_fd_sc_hd__o221a_2
XFILLER_156_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12023_ _13935_/Q vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13974_ _14095_/CLK _13974_/D vssd1 vssd1 vccd1 vccd1 _13974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ _12543_/X _12924_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12856_ _12525_/X input360/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _14398_/Q vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__inv_2
XPHY_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _09528_/X _12786_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13217_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14526_ _14527_/CLK _14526_/D vssd1 vssd1 vccd1 vccd1 _14526_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11738_ _11733_/Y _11689_/X _11734_/Y _11691_/X _11737_/X vssd1 vssd1 vccd1 vccd1
+ _11739_/D sky130_fd_sc_hd__o221a_1
XFILLER_109_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14457_ _14459_/CLK _14457_/D vssd1 vssd1 vccd1 vccd1 _14457_/Q sky130_fd_sc_hd__dfxtp_2
X_11669_ _11669_/A vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13408_ _14183_/CLK _13408_/D vssd1 vssd1 vccd1 vccd1 _13408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14388_ _14495_/CLK _14388_/D vssd1 vssd1 vccd1 vccd1 _14388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13339_ _13372_/CLK _13339_/D vssd1 vssd1 vccd1 vccd1 _13339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07900_ _14122_/Q _07892_/X _07726_/X _07894_/X _07897_/X vssd1 vssd1 vccd1 vccd1
+ _14122_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08880_ _08923_/A vssd1 vssd1 vccd1 vccd1 _08880_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07831_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07831_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07762_ _08153_/A vssd1 vssd1 vccd1 vccd1 _07762_/X sky130_fd_sc_hd__buf_4
XFILLER_110_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09501_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__clkbuf_2
X_06713_ _08822_/A vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07693_ _14214_/Q _07687_/X _07394_/X _07688_/X _07692_/X vssd1 vssd1 vccd1 vccd1
+ _14214_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ _09432_/A _12999_/X vssd1 vssd1 vccd1 vccd1 _13308_/D sky130_fd_sc_hd__and2_1
X_06644_ _06567_/Y input97/X _06696_/A _06588_/Y vssd1 vssd1 vccd1 vccd1 _06644_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09363_ _09364_/A _12839_/X vssd1 vssd1 vccd1 vccd1 _13364_/D sky130_fd_sc_hd__and2_1
X_06575_ input92/X vssd1 vssd1 vccd1 vccd1 _06575_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08314_ _13914_/Q _08310_/X _08153_/X _08311_/X _08313_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/D sky130_fd_sc_hd__o221a_1
X_09294_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_10 _11271_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _12030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_32 _08243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _13950_/Q _08237_/X _08158_/X _08238_/X _08239_/X vssd1 vssd1 vccd1 vccd1
+ _13950_/D sky130_fd_sc_hd__o221a_1
XANTENNA_43 _07370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_54 _07764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_65 _07929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_76 _08171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_87 _08632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _08176_/A vssd1 vssd1 vccd1 vccd1 _08176_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_98 _11660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07127_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07058_ _08243_/A vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__buf_4
XFILLER_118_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ _10962_/Y _10963_/X _10964_/Y _10965_/X _10970_/X vssd1 vssd1 vccd1 vccd1
+ _10992_/B sky130_fd_sc_hd__o221a_4
XFILLER_95_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12710_ _09565_/X _12709_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13690_ _14056_/CLK _13690_/D vssd1 vssd1 vccd1 vccd1 _13690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12641_ _13340_/Q _12640_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _13295_/Q _12571_/X input39/X vssd1 vssd1 vccd1 vccd1 _12572_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ _14527_/CLK _14311_/D vssd1 vssd1 vccd1 vccd1 _14311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _11521_/Y _11419_/X _11522_/Y _11421_/X vssd1 vssd1 vccd1 vccd1 _11523_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14242_ _14633_/CLK _14242_/D vssd1 vssd1 vccd1 vccd1 _14242_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11454_ _13922_/Q vssd1 vssd1 vccd1 vccd1 _11454_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10405_ _14603_/Q vssd1 vssd1 vccd1 vccd1 _10405_/Y sky130_fd_sc_hd__inv_2
X_14173_ _14173_/CLK _14173_/D vssd1 vssd1 vccd1 vccd1 _14173_/Q sky130_fd_sc_hd__dfxtp_1
X_11385_ _14272_/Q vssd1 vssd1 vccd1 vccd1 _11385_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _12641_/X input343/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__mux2_1
X_10336_ _14445_/Q vssd1 vssd1 vccd1 vccd1 _10336_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10267_ _10265_/Y _10181_/X _10266_/Y _10184_/X vssd1 vssd1 vccd1 vccd1 _10267_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13055_ _12606_/X _13054_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13055_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12006_ _13538_/Q vssd1 vssd1 vccd1 vccd1 _12006_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10198_ _10198_/A vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13957_ _13996_/CLK _13957_/D vssd1 vssd1 vccd1 vccd1 _13957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12908_ _12538_/X input349/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12908_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13888_ _14100_/CLK _13888_/D vssd1 vssd1 vccd1 vccd1 _13888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12839_ _12520_/X _12838_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12839_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ _14627_/CLK _14509_/D vssd1 vssd1 vccd1 vccd1 _14509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08030_ _14050_/Q _08025_/X _07710_/X _08027_/X _08017_/X vssd1 vssd1 vccd1 vccd1
+ _14050_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput30 io_in[36] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput41 la_data_in[101] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
XFILLER_156_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 la_data_in[111] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_1
XFILLER_11_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 la_data_in[121] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_1
XFILLER_176_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput74 la_data_in[16] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_1
XFILLER_143_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput85 la_data_in[26] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_1
Xinput96 la_data_in[36] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_4
XFILLER_196_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09981_ _09981_/A vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__inv_2
XFILLER_176_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08932_ _13601_/Q _08929_/X _08930_/X _08931_/X _08923_/X vssd1 vssd1 vccd1 vccd1
+ _13601_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08863_ _08871_/A vssd1 vssd1 vccd1 vccd1 _08863_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater620 _12858_/S vssd1 vssd1 vccd1 vccd1 _12922_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_84_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07814_ _14168_/Q _07808_/X _07708_/X _07811_/X _07812_/X vssd1 vssd1 vccd1 vccd1
+ _14168_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater631 _10076_/A vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__buf_6
XPHY_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater642 _14305_/CLK vssd1 vssd1 vccd1 vccd1 _14459_/CLK sky130_fd_sc_hd__clkbuf_8
XPHY_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater653 _14291_/CLK vssd1 vssd1 vccd1 vccd1 _14481_/CLK sky130_fd_sc_hd__buf_12
X_08794_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08794_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater664 _14123_/CLK vssd1 vssd1 vccd1 vccd1 _14094_/CLK sky130_fd_sc_hd__buf_12
XFILLER_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater675 _14110_/CLK vssd1 vssd1 vccd1 vccd1 _14107_/CLK sky130_fd_sc_hd__buf_12
XPHY_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater686 input78/X vssd1 vssd1 vccd1 vccd1 _12396_/S sky130_fd_sc_hd__buf_8
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07745_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07745_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater697 _13157_/S vssd1 vssd1 vccd1 vccd1 _13121_/S sky130_fd_sc_hd__buf_8
XPHY_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07676_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _09419_/A _13071_/X vssd1 vssd1 vccd1 vccd1 _13322_/D sky130_fd_sc_hd__and2_1
XFILLER_164_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06627_ _06545_/Y _06625_/Y _06545_/A _08920_/A vssd1 vssd1 vccd1 vccd1 _06627_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09346_ _09352_/A vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__clkbuf_2
X_06558_ _06558_/A vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09277_ _09277_/A vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__clkbuf_2
X_06489_ _09512_/A vssd1 vssd1 vccd1 vccd1 _13099_/S sky130_fd_sc_hd__clkinv_8
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08228_ _13960_/Q _08221_/X _08132_/X _08222_/X _08223_/X vssd1 vssd1 vccd1 vccd1
+ _13960_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08159_ _08184_/A vssd1 vssd1 vccd1 vccd1 _08159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11170_ _11406_/A vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10121_ _10126_/A _12454_/X vssd1 vssd1 vccd1 vccd1 _10121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10052_ _10052_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _10052_/Y sky130_fd_sc_hd__nor2_1
XPHY_7433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13811_ _14123_/CLK _13811_/D vssd1 vssd1 vccd1 vccd1 _13811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _14130_/CLK _13742_/D vssd1 vssd1 vccd1 vccd1 _13742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _11426_/A vssd1 vssd1 vccd1 vccd1 _10954_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13673_ _14071_/CLK _13673_/D vssd1 vssd1 vccd1 vccd1 _13673_/Q sky130_fd_sc_hd__dfxtp_1
X_10885_ _10883_/Y _10691_/X _10884_/Y _10693_/X vssd1 vssd1 vccd1 vccd1 _10885_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12624_ _09842_/X _13332_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12624_/X sky130_fd_sc_hd__mux2_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _13288_/Q _12554_/X _12619_/S vssd1 vssd1 vccd1 vccd1 _12555_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11487_/X _11506_/B _11506_/C _11506_/D vssd1 vssd1 vccd1 vccd1 _11507_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12486_ _12485_/X _06967_/Y _12486_/S vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14225_ _14459_/CLK _14225_/D vssd1 vssd1 vccd1 vccd1 _14225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11437_ _11437_/A vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14156_ _14305_/CLK _14156_/D vssd1 vssd1 vccd1 vccd1 _14156_/Q sky130_fd_sc_hd__dfxtp_1
X_11368_ _14116_/Q vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13107_ _12631_/X _13106_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
X_10319_ _13541_/Q _10206_/X _13782_/Q _10209_/X vssd1 vssd1 vccd1 vccd1 _10319_/X
+ sky130_fd_sc_hd__a22o_1
X_14087_ _14169_/CLK _14087_/D vssd1 vssd1 vccd1 vccd1 _14087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11299_ _11294_/Y _11199_/X _11295_/Y _11201_/X _11298_/X vssd1 vssd1 vccd1 vccd1
+ _11312_/B sky130_fd_sc_hd__o221a_1
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13038_ _13037_/X _12598_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07530_ _14302_/Q _07524_/X _07456_/X _07525_/X _07527_/X vssd1 vssd1 vccd1 vccd1
+ _14302_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07461_ _07476_/A vssd1 vssd1 vccd1 vccd1 _07461_/X sky130_fd_sc_hd__buf_1
XFILLER_126_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09200_ _13461_/Q _09135_/A _09060_/X _09137_/A _09196_/X vssd1 vssd1 vccd1 vccd1
+ _13461_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07392_ _08179_/A vssd1 vssd1 vccd1 vccd1 _07392_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09131_ _09131_/A _09271_/B _09131_/C _09271_/D vssd1 vssd1 vccd1 vccd1 _11693_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_143_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ _13539_/Q _08993_/A _09060_/X _08995_/A _09061_/X vssd1 vssd1 vccd1 vccd1
+ _13539_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _14058_/Q _08007_/X _07790_/X _08008_/X _08011_/X vssd1 vssd1 vccd1 vccd1
+ _14058_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09964_ _09888_/A _09888_/B _09889_/B vssd1 vssd1 vccd1 vccd1 _09964_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _13607_/Q _08905_/X _08914_/X _08907_/X _08910_/X vssd1 vssd1 vccd1 vccd1
+ _13607_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09895_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__or2_1
XFILLER_28_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08846_ _13645_/Q _08844_/X _08514_/X _08845_/X _08839_/X vssd1 vssd1 vccd1 vccd1
+ _13645_/D sky130_fd_sc_hd__o221a_1
XFILLER_150_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08777_ _08777_/A vssd1 vssd1 vccd1 vccd1 _08777_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07728_ _08119_/A vssd1 vssd1 vccd1 vccd1 _07728_/X sky130_fd_sc_hd__buf_4
XPHY_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07659_ _14234_/Q _07653_/X _07343_/X _07654_/X _07658_/X vssd1 vssd1 vccd1 vccd1
+ _14234_/D sky130_fd_sc_hd__o221a_1
XPHY_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10670_ _10668_/Y _10484_/X _10669_/Y _10487_/X vssd1 vssd1 vccd1 vccd1 _10670_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09329_ _13390_/Q _09326_/X _09051_/X _09327_/X _09322_/X vssd1 vssd1 vccd1 vccd1
+ _13390_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _12339_/X _13193_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12340_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12271_ _12061_/Y _13372_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12271_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14010_ _14130_/CLK _14010_/D vssd1 vssd1 vccd1 vccd1 _14010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _13481_/Q vssd1 vssd1 vccd1 vccd1 _11222_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ _14150_/Q vssd1 vssd1 vccd1 vccd1 _11153_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10138_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__buf_1
XFILLER_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11084_ _13401_/Q _11042_/X _13713_/Q _10936_/X vssd1 vssd1 vccd1 vccd1 _11084_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_7230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput220 la_oenb[32] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_1
XPHY_7241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput231 la_oenb[42] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_1
XPHY_7252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _13372_/Q _10002_/B _10003_/A vssd1 vssd1 vccd1 vccd1 _10035_/X sky130_fd_sc_hd__o21a_1
Xinput242 la_oenb[52] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_1
XFILLER_81_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput253 la_oenb[62] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__buf_1
XFILLER_23_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput264 la_oenb[72] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_hd__buf_1
XPHY_7285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput275 la_oenb[82] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_hd__buf_1
XPHY_7296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput286 la_oenb[92] vssd1 vssd1 vccd1 vccd1 input286/X sky130_fd_sc_hd__buf_1
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput297 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _06499_/B sky130_fd_sc_hd__buf_1
XPHY_6573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _11984_/Y _10248_/A _11985_/Y _10251_/A vssd1 vssd1 vccd1 vccd1 _11986_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13725_ _14178_/CLK _13725_/D vssd1 vssd1 vccd1 vccd1 _13725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10937_ _13398_/Q _10804_/X _13710_/Q _10936_/X vssd1 vssd1 vccd1 vccd1 _10937_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13656_ _14056_/CLK _13656_/D vssd1 vssd1 vccd1 vccd1 _13656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10868_ _13591_/Q vssd1 vssd1 vccd1 vccd1 _10868_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _09855_/X _13325_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__mux2_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13587_ _14183_/CLK _13587_/D vssd1 vssd1 vccd1 vccd1 _13587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ _13434_/Q vssd1 vssd1 vccd1 vccd1 _10799_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12538_ _13378_/Q _10018_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12469_ _12468_/X _06943_/X _12502_/S vssd1 vssd1 vccd1 vccd1 _12469_/X sky130_fd_sc_hd__mux2_2
X_14208_ _14325_/CLK _14208_/D vssd1 vssd1 vccd1 vccd1 _14208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ _14139_/CLK _14139_/D vssd1 vssd1 vccd1 vccd1 _14139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06961_ _14572_/Q vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08700_ _13723_/Q _08698_/X _08514_/X _08699_/X _08696_/X vssd1 vssd1 vccd1 vccd1
+ _13723_/D sky130_fd_sc_hd__o221a_1
XFILLER_45_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09680_ _09726_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__or2_1
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06892_ _14590_/Q vssd1 vssd1 vccd1 vccd1 _06893_/A sky130_fd_sc_hd__inv_2
XFILLER_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08631_ _13757_/Q _08626_/X _08546_/X _08627_/X _08628_/X vssd1 vssd1 vccd1 vccd1
+ _13757_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08562_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08562_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07513_ _14313_/Q _07508_/X _07341_/X _07509_/X _07511_/X vssd1 vssd1 vccd1 vccd1
+ _14313_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08493_ _13816_/Q _08486_/X _08492_/X _08488_/X _08480_/X vssd1 vssd1 vccd1 vccd1
+ _13816_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07444_ _07476_/A vssd1 vssd1 vccd1 vccd1 _07444_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07375_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _13512_/Q _09111_/X _08960_/X _09112_/X _09109_/X vssd1 vssd1 vccd1 vccd1
+ _13512_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09045_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09947_ _09891_/A _09891_/B _09946_/Y vssd1 vssd1 vccd1 vccd1 _09947_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09878_ _13290_/Q vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__inv_2
XFILLER_63_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08829_ _08829_/A vssd1 vssd1 vccd1 vccd1 _08829_/X sky130_fd_sc_hd__buf_4
XPHY_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11840_ _11838_/Y _11653_/X _11839_/Y _11655_/X vssd1 vssd1 vccd1 vccd1 _11840_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11771_ _14202_/Q vssd1 vssd1 vccd1 vccd1 _11771_/Y sky130_fd_sc_hd__inv_2
XPHY_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13510_ _14110_/CLK _13510_/D vssd1 vssd1 vccd1 vccd1 _13510_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _13549_/Q _10720_/X _13790_/Q _10721_/X vssd1 vssd1 vccd1 vccd1 _10722_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14490_ _14611_/CLK _14490_/D vssd1 vssd1 vccd1 vccd1 _14490_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _14188_/CLK _13441_/D vssd1 vssd1 vccd1 vccd1 _13441_/Q sky130_fd_sc_hd__dfxtp_1
X_10653_ _13945_/Q vssd1 vssd1 vccd1 vccd1 _10653_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ _13372_/CLK _13372_/D vssd1 vssd1 vccd1 vccd1 _13372_/Q sky130_fd_sc_hd__dfxtp_1
X_10584_ _14489_/Q vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _13198_/Q _06829_/Y _12368_/S vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ _12038_/Y _13355_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11205_ _11441_/A vssd1 vssd1 vccd1 vccd1 _11205_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12185_ vssd1 vssd1 vccd1 vccd1 _12185_/HI _12185_/LO sky130_fd_sc_hd__conb_1
XFILLER_46_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11136_ _11134_/Y _10952_/X _11135_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _11136_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11067_ _14265_/Q vssd1 vssd1 vccd1 vccd1 _11067_/Y sky130_fd_sc_hd__inv_2
XPHY_7060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _13378_/Q _10017_/B _10019_/A vssd1 vssd1 vccd1 vccd1 _10018_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11969_ _13732_/Q _10173_/A _14051_/Q _10203_/A _11968_/X vssd1 vssd1 vccd1 vccd1
+ _11969_/X sky130_fd_sc_hd__a221o_2
XFILLER_127_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13708_ _14183_/CLK _13708_/D vssd1 vssd1 vccd1 vccd1 _13708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13639_ _14146_/CLK _13639_/D vssd1 vssd1 vccd1 vccd1 _13639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07160_ _08744_/A _09063_/B _09271_/C _09271_/D vssd1 vssd1 vccd1 vccd1 _11695_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_53_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07091_ _07144_/A vssd1 vssd1 vccd1 vccd1 _07092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput502 _12133_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__clkbuf_2
Xoutput513 _12143_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__clkbuf_2
Xoutput524 _12153_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput535 _12163_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput546 _12173_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__clkbuf_2
Xoutput557 _12183_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput568 _12193_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput579 _13267_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _09801_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__or2_1
XFILLER_64_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07993_ _14071_/Q _07991_/X _07759_/X _07992_/X _07987_/X vssd1 vssd1 vccd1 vccd1
+ _14071_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _09732_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__and2_1
XFILLER_5_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06944_ _06937_/X _12305_/X _06943_/X _06939_/X vssd1 vssd1 vccd1 vccd1 _06945_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09663_ _09732_/A _10070_/A vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__nand2_4
XFILLER_3_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06875_ _14594_/Q vssd1 vssd1 vccd1 vccd1 _06875_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08614_ _13768_/Q _08610_/X _08517_/X _08611_/X _08612_/X vssd1 vssd1 vccd1 vccd1
+ _13768_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _09583_/X _09593_/X _13257_/Q _09584_/X vssd1 vssd1 vccd1 vccd1 _13225_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _13797_/Q _08540_/X _08544_/X _08542_/X _08538_/X vssd1 vssd1 vccd1 vccd1
+ _13797_/D sky130_fd_sc_hd__o221a_1
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08476_ _13823_/Q _08468_/X _08183_/X _08469_/X _08474_/X vssd1 vssd1 vccd1 vccd1
+ _13823_/D sky130_fd_sc_hd__o221a_1
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07427_ _14358_/Q _07422_/X _07327_/X _07424_/X _07425_/X vssd1 vssd1 vccd1 vccd1
+ _14358_/D sky130_fd_sc_hd__o221a_1
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _08146_/A vssd1 vssd1 vccd1 vccd1 _07358_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07289_ _14413_/Q _07282_/X _06820_/X _07283_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _14413_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09028_ _13559_/Q _09022_/X _08940_/X _09023_/X _09027_/X vssd1 vssd1 vccd1 vccd1
+ _13559_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13990_ _14107_/CLK _13990_/D vssd1 vssd1 vccd1 vccd1 _13990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12941_ _12551_/X _12940_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12872_ _12529_/X input342/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__mux2_1
XANTENNA_100 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_111 _11451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/CLK _14611_/D vssd1 vssd1 vccd1 vccd1 _14611_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_122 _10838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ _11823_/A _11823_/B _11823_/C _11823_/D vssd1 vssd1 vccd1 vccd1 _11823_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_155 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_177 input333/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ _14621_/CLK _14542_/D vssd1 vssd1 vccd1 vccd1 _14542_/Q sky130_fd_sc_hd__dfxtp_1
X_11754_ _13851_/Q vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 input351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 input361/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10705_ _13868_/Q vssd1 vssd1 vccd1 vccd1 _10705_/Y sky130_fd_sc_hd__inv_2
XPHY_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14473_ _14527_/CLK _14473_/D vssd1 vssd1 vccd1 vccd1 _14473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _11685_/A vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__buf_2
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13424_ _14056_/CLK _13424_/D vssd1 vssd1 vccd1 vccd1 _13424_/Q sky130_fd_sc_hd__dfxtp_1
X_10636_ _10631_/Y _10492_/X _10632_/Y _10495_/X _10635_/X vssd1 vssd1 vccd1 vccd1
+ _10643_/C sky130_fd_sc_hd__o221a_1
XFILLER_161_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13355_ _14639_/CLK _13355_/D vssd1 vssd1 vccd1 vccd1 _13355_/Q sky130_fd_sc_hd__dfxtp_1
X_10567_ _10562_/Y _10425_/X _10563_/Y _10428_/X _10566_/X vssd1 vssd1 vccd1 vccd1
+ _10603_/A sky130_fd_sc_hd__o221a_2
XFILLER_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12306_ _11035_/Y _14537_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12306_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13286_ _14538_/CLK _13286_/D vssd1 vssd1 vccd1 vccd1 _13286_/Q sky130_fd_sc_hd__dfxtp_4
X_10498_ _11449_/A vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12237_ _12237_/A vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12168_ vssd1 vssd1 vccd1 vccd1 _12168_/HI _12168_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11119_ _14072_/Q vssd1 vssd1 vccd1 vccd1 _11119_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ vssd1 vssd1 vccd1 vccd1 _12099_/HI _12099_/LO sky130_fd_sc_hd__conb_1
XFILLER_81_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XFILLER_42_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06660_ _06567_/Y _06659_/X _06567_/Y _06659_/X vssd1 vssd1 vccd1 vccd1 _06660_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06591_ input95/X vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08330_ _13904_/Q _08326_/X _08259_/X _08327_/X _08329_/X vssd1 vssd1 vccd1 vccd1
+ _13904_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08261_ _13942_/Q _08255_/X _08179_/X _08256_/X _08257_/X vssd1 vssd1 vccd1 vccd1
+ _13942_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07212_ _14455_/Q _07209_/X _06810_/X _07210_/X _07205_/X vssd1 vssd1 vccd1 vccd1
+ _14455_/D sky130_fd_sc_hd__o221a_1
XFILLER_18_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08192_ _13975_/Q _08095_/A _07876_/X _08097_/A _08184_/X vssd1 vssd1 vccd1 vccd1
+ _13975_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07143_ _14491_/Q _07136_/X _06820_/X _07137_/X _07139_/X vssd1 vssd1 vccd1 vccd1
+ _14491_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07074_ _14528_/Q _07069_/X _07073_/X _07070_/X _07071_/X vssd1 vssd1 vccd1 vccd1
+ _14528_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput376 _12213_/X vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput387 _12223_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput398 _12075_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07976_ _14081_/Q _07974_/X _07733_/X _07975_/X _07970_/X vssd1 vssd1 vccd1 vccd1
+ _14081_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _06943_/X _09702_/X _06943_/X _09702_/X vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06927_ _14581_/Q vssd1 vssd1 vccd1 vccd1 _06927_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09646_ _09637_/Y _09645_/X _09637_/Y _09645_/X vssd1 vssd1 vccd1 vccd1 _09646_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06858_ _14598_/Q vssd1 vssd1 vccd1 vccd1 _06858_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09577_ _09570_/X _09576_/X _13264_/Q _09571_/X vssd1 vssd1 vccd1 vccd1 _13232_/D
+ sky130_fd_sc_hd__o22a_1
X_06789_ _08150_/A vssd1 vssd1 vccd1 vccd1 _06789_/X sky130_fd_sc_hd__clkbuf_4
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08554_/A vssd1 vssd1 vccd1 vccd1 _08528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _13833_/Q _08452_/X _08158_/X _08453_/X _08457_/X vssd1 vssd1 vccd1 vccd1
+ _13833_/D sky130_fd_sc_hd__o221a_1
XFILLER_141_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11470_ _11468_/Y _11401_/X _11469_/Y _11403_/X vssd1 vssd1 vccd1 vccd1 _11470_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10402_/X _10421_/B _10421_/C _10421_/D vssd1 vssd1 vccd1 vccd1 _10422_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_123_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13140_ _12649_/X input338/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__mux2_1
X_10352_ _10350_/Y _10181_/X _10351_/Y _10184_/X vssd1 vssd1 vccd1 vccd1 _10352_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _12614_/X _13070_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13071_/X sky130_fd_sc_hd__mux2_1
X_10283_ _10281_/Y _10220_/X _10282_/Y _10223_/X vssd1 vssd1 vccd1 vccd1 _10283_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12022_ _12017_/Y _10228_/A _12018_/Y _10231_/A _12021_/X vssd1 vssd1 vccd1 vccd1
+ _12029_/C sky130_fd_sc_hd__o221a_1
XFILLER_152_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13973_ _14095_/CLK _13973_/D vssd1 vssd1 vccd1 vccd1 _13973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12924_ _12543_/X input359/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12855_ _12524_/X _12854_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _14632_/Q vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__inv_2
XPHY_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ _09528_/X _12785_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14525_ _14527_/CLK _14525_/D vssd1 vssd1 vccd1 vccd1 _14525_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11737_ _11735_/Y _11693_/X _11736_/Y _11695_/X vssd1 vssd1 vccd1 vccd1 _11737_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14470_/CLK _14456_/D vssd1 vssd1 vccd1 vccd1 _14456_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11668_ _14512_/Q vssd1 vssd1 vccd1 vccd1 _11668_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _14183_/CLK _13407_/D vssd1 vssd1 vccd1 vccd1 _13407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10619_ _13983_/Q vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__inv_2
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14387_ _14495_/CLK _14387_/D vssd1 vssd1 vccd1 vccd1 _14387_/Q sky130_fd_sc_hd__dfxtp_1
X_11599_ _13965_/Q vssd1 vssd1 vccd1 vccd1 _11599_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13338_ _13370_/CLK _13338_/D vssd1 vssd1 vccd1 vccd1 _13338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13269_ _14639_/CLK _13269_/D vssd1 vssd1 vccd1 vccd1 _13269_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07830_ _07856_/A vssd1 vssd1 vccd1 vccd1 _07830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07761_ _14188_/Q _07758_/X _07759_/X _07760_/X _07756_/X vssd1 vssd1 vccd1 vccd1
+ _14188_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09500_ _09500_/A vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__clkbuf_2
X_06712_ _14637_/Q _06530_/X _06532_/X _07809_/A _06723_/C1 vssd1 vssd1 vccd1 vccd1
+ _14637_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07692_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07692_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09431_ _09432_/A _12995_/X vssd1 vssd1 vccd1 vccd1 _13309_/D sky130_fd_sc_hd__and2_1
X_06643_ _06634_/X _06642_/X _06634_/X _06642_/X vssd1 vssd1 vccd1 vccd1 _06643_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09362_ _09364_/A _12835_/X vssd1 vssd1 vccd1 vccd1 _13365_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06574_ input94/X vssd1 vssd1 vccd1 vccd1 _06574_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08313_ _08329_/A vssd1 vssd1 vccd1 vccd1 _08313_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09293_ _13412_/Q _09285_/X _08119_/A _09287_/X _09290_/X vssd1 vssd1 vccd1 vccd1
+ _13412_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_11 _11313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _09732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08244_ _13951_/Q _08237_/X _08243_/X _08238_/X _08239_/X vssd1 vssd1 vccd1 vccd1
+ _13951_/D sky130_fd_sc_hd__o221a_1
XANTENNA_33 _08243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _07370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_55 _07767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 _07960_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_77 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_88 _08653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__buf_4
XFILLER_119_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_99 _09173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ _14501_/Q _07119_/X _06784_/X _07120_/X _07122_/X vssd1 vssd1 vccd1 vccd1
+ _14501_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07057_ _14537_/Q _07052_/X _06796_/X _07053_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _14537_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07959_ _14090_/Q _07955_/X _07708_/X _07957_/X _07946_/X vssd1 vssd1 vccd1 vccd1
+ _14090_/D sky130_fd_sc_hd__o221a_1
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10970_ _10966_/Y _10967_/X _10968_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _10970_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ _14594_/Q _14585_/Q _06875_/Y _06912_/Y vssd1 vssd1 vccd1 vccd1 _09629_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12640_ _09829_/X _13340_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__mux2_1
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12571_ _09944_/Y _13295_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _14495_/CLK _14310_/D vssd1 vssd1 vccd1 vccd1 _14310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11522_ _14119_/Q vssd1 vssd1 vccd1 vccd1 _11522_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14241_ _14633_/CLK _14241_/D vssd1 vssd1 vccd1 vccd1 _14241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _11444_/Y _11445_/X _11446_/Y _11447_/X _11452_/X vssd1 vssd1 vccd1 vccd1
+ _11464_/C sky130_fd_sc_hd__o221a_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10404_ _14330_/Q vssd1 vssd1 vccd1 vccd1 _10404_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14172_ _14173_/CLK _14172_/D vssd1 vssd1 vccd1 vccd1 _14172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11384_ _14194_/Q vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13123_ _12639_/X _13122_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ _13463_/Q vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13054_ _13053_/X _12606_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13054_/X sky130_fd_sc_hd__mux2_1
X_10266_ _13859_/Q vssd1 vssd1 vccd1 vccd1 _10266_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12005_ _14013_/Q vssd1 vssd1 vccd1 vccd1 _12005_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10197_ _11660_/A vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__buf_2
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13956_ _13996_/CLK _13956_/D vssd1 vssd1 vccd1 vccd1 _13956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _12537_/X _12906_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13887_ _14100_/CLK _13887_/D vssd1 vssd1 vccd1 vccd1 _13887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12838_ _12520_/X _12837_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12769_ _09519_/X _12768_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14508_ _14627_/CLK _14508_/D vssd1 vssd1 vccd1 vccd1 _14508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 io_in[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
Xinput31 io_in[37] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
X_14439_ _14481_/CLK _14439_/D vssd1 vssd1 vccd1 vccd1 _14439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 la_data_in[102] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
Xinput53 la_data_in[112] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_1
Xinput64 la_data_in[122] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
XFILLER_7_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput75 la_data_in[17] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 la_data_in[27] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
XFILLER_176_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 la_data_in[37] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__buf_2
XFILLER_196_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09980_ _13361_/Q _09980_/B vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08931_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08931_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _13635_/Q _08860_/X _08541_/X _08861_/X _08855_/X vssd1 vssd1 vccd1 vccd1
+ _13635_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater610 _12666_/S vssd1 vssd1 vccd1 vccd1 _12658_/S sky130_fd_sc_hd__buf_6
X_07813_ _14169_/Q _07808_/X _07809_/X _07811_/X _07812_/X vssd1 vssd1 vccd1 vccd1
+ _14169_/D sky130_fd_sc_hd__o221a_1
Xrepeater621 _12407_/S vssd1 vssd1 vccd1 vccd1 _12416_/S sky130_fd_sc_hd__buf_8
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _08793_/A vssd1 vssd1 vccd1 vccd1 _08793_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater632 _06918_/A vssd1 vssd1 vccd1 vccd1 _06515_/A1 sky130_fd_sc_hd__buf_6
XPHY_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater643 _14470_/CLK vssd1 vssd1 vccd1 vccd1 _14305_/CLK sky130_fd_sc_hd__buf_12
XFILLER_211_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater654 _14529_/CLK vssd1 vssd1 vccd1 vccd1 _14291_/CLK sky130_fd_sc_hd__buf_6
XFILLER_113_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater665 _14121_/CLK vssd1 vssd1 vccd1 vccd1 _14123_/CLK sky130_fd_sc_hd__buf_6
XFILLER_42_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07744_ _14194_/Q _07732_/X _07742_/X _07734_/X _07743_/X vssd1 vssd1 vccd1 vccd1
+ _14194_/D sky130_fd_sc_hd__o221a_1
Xrepeater676 _13996_/CLK vssd1 vssd1 vccd1 vccd1 _14110_/CLK sky130_fd_sc_hd__buf_12
XPHY_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater687 _12659_/S vssd1 vssd1 vccd1 vccd1 _12667_/S sky130_fd_sc_hd__buf_8
Xrepeater698 _13133_/S vssd1 vssd1 vccd1 vccd1 _13157_/S sky130_fd_sc_hd__buf_8
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07675_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__buf_2
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09414_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__buf_4
XFILLER_198_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06626_ _06626_/A vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09345_ _09345_/A _12911_/X vssd1 vssd1 vccd1 vccd1 _13378_/D sky130_fd_sc_hd__and2_1
XFILLER_107_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ _06559_/A vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__buf_2
XFILLER_70_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09276_ _09327_/A vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06488_ _06488_/A _06488_/B vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__nand2_8
XFILLER_33_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08227_ _13961_/Q _08221_/X _08130_/X _08222_/X _08223_/X vssd1 vssd1 vccd1 vccd1
+ _13961_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _08158_/A vssd1 vssd1 vccd1 vccd1 _08158_/X sky130_fd_sc_hd__buf_4
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07109_ _14512_/Q _07102_/X _06745_/X _07104_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _14512_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08089_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08089_/X sky130_fd_sc_hd__buf_2
XFILLER_106_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _12452_/S sky130_fd_sc_hd__or2_1
XFILLER_134_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ _13353_/Q _09967_/B _13354_/Q vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__a21oi_1
XPHY_7423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13810_ _14123_/CLK _13810_/D vssd1 vssd1 vccd1 vccd1 _13810_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_6777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13741_ _14130_/CLK _13741_/D vssd1 vssd1 vccd1 vccd1 _13741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10953_ _13515_/Q vssd1 vssd1 vccd1 vccd1 _10953_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13672_ _14071_/CLK _13672_/D vssd1 vssd1 vccd1 vccd1 _13672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10884_ _13631_/Q vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ _13333_/Q _12622_/X input39/X vssd1 vssd1 vccd1 vccd1 _12623_/X sky130_fd_sc_hd__mux2_1
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _09956_/X _13288_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11500_/Y _11455_/X _11501_/Y _11457_/X _11504_/X vssd1 vssd1 vccd1 vccd1
+ _11506_/D sky130_fd_sc_hd__o221a_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ _12509_/X _06967_/Y _12485_/S vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14224_ _14459_/CLK _14224_/D vssd1 vssd1 vccd1 vccd1 _14224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11436_ _14351_/Q vssd1 vssd1 vccd1 vccd1 _11436_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14155_ _14470_/CLK _14155_/D vssd1 vssd1 vccd1 vccd1 _14155_/Q sky130_fd_sc_hd__dfxtp_1
X_11367_ _13843_/Q vssd1 vssd1 vccd1 vccd1 _11367_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _13105_/X _12631_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__mux2_1
X_10318_ _10308_/Y _10178_/X _10311_/X _10314_/X _10317_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/C sky130_fd_sc_hd__o2111a_4
XFILLER_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14086_ _14178_/CLK _14086_/D vssd1 vssd1 vccd1 vccd1 _14086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11298_ _11296_/Y _11203_/X _11297_/Y _11205_/X vssd1 vssd1 vccd1 vccd1 _11298_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13037_ _12598_/X _13036_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10249_ _14443_/Q vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _14095_/CLK _13939_/D vssd1 vssd1 vccd1 vccd1 _13939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07460_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07391_ _14372_/Q _07387_/X _07073_/X _07389_/X _07385_/X vssd1 vssd1 vccd1 vccd1
+ _14372_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09130_ _13500_/Q _09067_/A _09060_/X _09069_/A _09125_/X vssd1 vssd1 vccd1 vccd1
+ _13500_/D sky130_fd_sc_hd__o221a_1
XFILLER_56_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09061_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09061_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08012_ _14059_/Q _08007_/X _07788_/X _08008_/X _08011_/X vssd1 vssd1 vccd1 vccd1
+ _14059_/D sky130_fd_sc_hd__o221a_1
XFILLER_89_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09963_ _13293_/Q _09961_/Y _09888_/B vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08914_ _08914_/A vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__buf_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09894_ _09894_/A _09949_/A vssd1 vssd1 vccd1 vccd1 _09895_/B sky130_fd_sc_hd__or2_1
XFILLER_24_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08869_/A vssd1 vssd1 vccd1 vccd1 _08845_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08776_ _08793_/A vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07727_ _14200_/Q _07718_/X _07726_/X _07721_/X _07715_/X vssd1 vssd1 vccd1 vccd1
+ _14200_/D sky130_fd_sc_hd__o221a_1
XPHY_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07658_/X sky130_fd_sc_hd__buf_2
XPHY_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06609_ _06609_/A vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_198_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07589_ _07605_/A vssd1 vssd1 vccd1 vccd1 _07589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09328_ _13391_/Q _09326_/X _08175_/A _09327_/X _09322_/X vssd1 vssd1 vccd1 vccd1
+ _13391_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09259_ _13430_/Q _09257_/X _08970_/X _09258_/X _09252_/X vssd1 vssd1 vccd1 vccd1
+ _13430_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12270_ _12060_/Y _13371_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11221_ _11457_/A vssd1 vssd1 vccd1 vccd1 _11221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11152_ _13916_/Q vssd1 vssd1 vccd1 vccd1 _11152_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ _12508_/S _10103_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__or2_2
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11083_ _11078_/Y _10923_/X _11079_/Y _10925_/X _11082_/X vssd1 vssd1 vccd1 vccd1
+ _11118_/A sky130_fd_sc_hd__o221a_2
XPHY_7220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput210 la_oenb[23] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__buf_1
XFILLER_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput221 la_oenb[33] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_1
X_10034_ _13371_/Q _10000_/B _10001_/A vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__o21a_1
Xinput232 la_oenb[43] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_1
XPHY_7253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 la_oenb[53] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_1
XFILLER_209_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput254 la_oenb[63] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__buf_1
XFILLER_76_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput265 la_oenb[73] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_hd__buf_1
XFILLER_40_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput276 la_oenb[83] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_hd__buf_1
XPHY_7297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput287 la_oenb[93] vssd1 vssd1 vccd1 vccd1 input287/X sky130_fd_sc_hd__buf_1
XPHY_6563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput298 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _06503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _14480_/Q vssd1 vssd1 vccd1 vccd1 _11985_/Y sky130_fd_sc_hd__inv_2
XPHY_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13724_ _14178_/CLK _13724_/D vssd1 vssd1 vccd1 vccd1 _13724_/Q sky130_fd_sc_hd__dfxtp_1
X_10936_ _11408_/A vssd1 vssd1 vccd1 vccd1 _10936_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13655_ _14056_/CLK _13655_/D vssd1 vssd1 vccd1 vccd1 _13655_/Q sky130_fd_sc_hd__dfxtp_1
X_10867_ _14300_/Q vssd1 vssd1 vccd1 vccd1 _10867_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _13326_/Q _12605_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12606_/X sky130_fd_sc_hd__mux2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _14178_/CLK _13586_/D vssd1 vssd1 vccd1 vccd1 _13586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _14065_/Q vssd1 vssd1 vccd1 vccd1 _10798_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12537_ _13379_/Q _10021_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12537_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12467_/X _06943_/X _12603_/S vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14207_ _14325_/CLK _14207_/D vssd1 vssd1 vccd1 vccd1 _14207_/Q sky130_fd_sc_hd__dfxtp_1
X_11419_ _11419_/A vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12399_ _13221_/Q _12398_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14138_ _14139_/CLK _14138_/D vssd1 vssd1 vccd1 vccd1 _14138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06960_ _06972_/A _06960_/B vssd1 vssd1 vccd1 vccd1 _14573_/D sky130_fd_sc_hd__nor2_1
X_14069_ _14071_/CLK _14069_/D vssd1 vssd1 vccd1 vccd1 _14069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06891_ _06899_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _14591_/D sky130_fd_sc_hd__nor2_1
X_08630_ _13758_/Q _08626_/X _08544_/X _08627_/X _08628_/X vssd1 vssd1 vccd1 vccd1
+ _13758_/D sky130_fd_sc_hd__o221a_1
XFILLER_23_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08561_ _13790_/Q _08552_/X _08560_/X _08554_/X _08550_/X vssd1 vssd1 vccd1 vccd1
+ _13790_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07512_ _14314_/Q _07508_/X _07339_/X _07509_/X _07511_/X vssd1 vssd1 vccd1 vccd1
+ _14314_/D sky130_fd_sc_hd__o221a_1
XFILLER_184_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _08825_/A vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__buf_2
XFILLER_1_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07374_ _08162_/A vssd1 vssd1 vccd1 vccd1 _07374_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_206_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09113_ _13513_/Q _09111_/X _08957_/X _09112_/X _09109_/X vssd1 vssd1 vccd1 vccd1
+ _13513_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09044_ _09138_/A vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__buf_2
XFILLER_191_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09946_ _09946_/A vssd1 vssd1 vccd1 vccd1 _09946_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09877_ _13291_/Q vssd1 vssd1 vccd1 vccd1 _09885_/A sky130_fd_sc_hd__inv_2
XFILLER_189_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08828_ _13652_/Q _08818_/X _08827_/X _08820_/X _08823_/X vssd1 vssd1 vccd1 vccd1
+ _13652_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08801_/A vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__buf_4
XFILLER_76_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _13610_/Q vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__inv_2
XPHY_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10721_ _11431_/A vssd1 vssd1 vccd1 vccd1 _10721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13440_ _14146_/CLK _13440_/D vssd1 vssd1 vccd1 vccd1 _13440_/Q sky130_fd_sc_hd__dfxtp_1
X_10652_ _14218_/Q _10437_/X _14413_/Q _10438_/X _10651_/X vssd1 vssd1 vccd1 vccd1
+ _10685_/B sky130_fd_sc_hd__a221oi_2
XFILLER_74_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13371_ _13371_/CLK _13371_/D vssd1 vssd1 vccd1 vccd1 _13371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10583_ _13198_/Q _10539_/X _14021_/Q _10469_/X _10582_/X vssd1 vssd1 vccd1 vccd1
+ _10583_/X sky130_fd_sc_hd__a221o_4
XFILLER_107_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12322_ _10255_/Y _14521_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12322_/X sky130_fd_sc_hd__mux2_4
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12253_ _12034_/Y _13354_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12253_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _14385_/Q vssd1 vssd1 vccd1 vccd1 _11204_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ vssd1 vssd1 vccd1 vccd1 _12184_/HI _12184_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11135_ _13519_/Q vssd1 vssd1 vccd1 vccd1 _11135_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11066_ _14187_/Q vssd1 vssd1 vccd1 vccd1 _11066_/Y sky130_fd_sc_hd__inv_2
XPHY_7050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _13378_/Q _10017_/B vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11968_ _13576_/Q _10206_/A _13817_/Q _10209_/A vssd1 vssd1 vccd1 vccd1 _11968_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ _14183_/CLK _13707_/D vssd1 vssd1 vccd1 vccd1 _13707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _10914_/Y _10745_/X _10915_/Y _10747_/X _10918_/X vssd1 vssd1 vccd1 vccd1
+ _10920_/D sky130_fd_sc_hd__o221a_1
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11899_ _11894_/Y _10228_/A _11895_/Y _10231_/A _11898_/X vssd1 vssd1 vccd1 vccd1
+ _11906_/C sky130_fd_sc_hd__o221a_1
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _14146_/CLK _13638_/D vssd1 vssd1 vccd1 vccd1 _13638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13569_ _14121_/CLK _13569_/D vssd1 vssd1 vccd1 vccd1 _13569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07090_ _07145_/A vssd1 vssd1 vccd1 vccd1 _07144_/A sky130_fd_sc_hd__inv_2
XFILLER_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput503 _12134_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput514 _12144_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput525 _12154_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput536 _12164_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput547 _12174_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__clkbuf_2
Xoutput558 _12184_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput569 _12194_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09800_ _13345_/Q vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__inv_2
XFILLER_64_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ _08000_/A vssd1 vssd1 vccd1 vccd1 _07992_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06943_ _06943_/A vssd1 vssd1 vccd1 vccd1 _06943_/X sky130_fd_sc_hd__clkbuf_4
X_09731_ _09727_/X _09730_/X _09727_/X _09730_/X vssd1 vssd1 vccd1 vccd1 _10103_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09662_ _09642_/X _09661_/X _09642_/X _09661_/X vssd1 vssd1 vccd1 vccd1 _10070_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_3_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06874_ _06877_/A _06874_/B vssd1 vssd1 vccd1 vccd1 _14595_/D sky130_fd_sc_hd__nor2_1
X_08613_ _13769_/Q _08610_/X _08514_/X _08611_/X _08612_/X vssd1 vssd1 vccd1 vccd1
+ _13769_/D sky130_fd_sc_hd__o221a_1
XFILLER_209_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09593_ _09597_/A _12340_/X vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__and2_1
XFILLER_209_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08544_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08544_/X sky130_fd_sc_hd__clkbuf_4
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _13824_/Q _08468_/X _08181_/X _08469_/X _08474_/X vssd1 vssd1 vccd1 vccd1
+ _13824_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07426_ _14359_/Q _07422_/X _07323_/X _07424_/X _07425_/X vssd1 vssd1 vccd1 vccd1
+ _14359_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07357_ _14385_/Q _07348_/X _07356_/X _07350_/X _07346_/X vssd1 vssd1 vccd1 vccd1
+ _14385_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07288_ _14414_/Q _07282_/X _06817_/X _07283_/X _07287_/X vssd1 vssd1 vccd1 vccd1
+ _14414_/D sky130_fd_sc_hd__o221a_1
X_09027_ _09036_/A vssd1 vssd1 vccd1 vccd1 _09027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09929_ _13318_/Q vssd1 vssd1 vccd1 vccd1 _09929_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12940_ _12551_/X input355/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12528_/X _12870_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12871_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_101 _09236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _11455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _14627_/CLK _14610_/D vssd1 vssd1 vccd1 vccd1 _14610_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_123 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ _11803_/X _11822_/B _11822_/C _11822_/D vssd1 vssd1 vccd1 vccd1 _11823_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_134 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_156 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_167 _12029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11753_ _11751_/Y _11648_/X _11752_/Y _11650_/X vssd1 vssd1 vccd1 vccd1 _11753_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_178 input333/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ _14621_/CLK _14541_/D vssd1 vssd1 vccd1 vccd1 _14541_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 input352/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11414_/A vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _14278_/Q vssd1 vssd1 vccd1 vccd1 _11684_/Y sky130_fd_sc_hd__inv_2
X_14472_ _14527_/CLK _14472_/D vssd1 vssd1 vccd1 vccd1 _14472_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _14056_/CLK _13423_/D vssd1 vssd1 vccd1 vccd1 _13423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10635_ _10633_/Y _10498_/X _10634_/Y _10501_/X vssd1 vssd1 vccd1 vccd1 _10635_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13354_ _14639_/CLK _13354_/D vssd1 vssd1 vccd1 vccd1 _13354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10566_ _10564_/Y _10431_/X _10565_/Y _10434_/X vssd1 vssd1 vccd1 vccd1 _10566_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _11077_/Y _14538_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12305_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13285_ _14538_/CLK _13285_/D vssd1 vssd1 vccd1 vccd1 _13285_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10497_ _11683_/A vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__buf_4
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _12236_/A vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12167_ vssd1 vssd1 vccd1 vccd1 _12167_/HI _12167_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11118_ _11118_/A _11118_/B _11118_/C _11118_/D vssd1 vssd1 vccd1 vccd1 _11118_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12098_ vssd1 vssd1 vccd1 vccd1 _12098_/HI _12098_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11049_ _13836_/Q vssd1 vssd1 vccd1 vccd1 _11049_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_42_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06590_ input97/X vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__buf_2
XFILLER_94_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08260_ _13943_/Q _08255_/X _08259_/X _08256_/X _08257_/X vssd1 vssd1 vccd1 vccd1
+ _13943_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ _14456_/Q _07209_/X _06807_/X _07210_/X _07205_/X vssd1 vssd1 vccd1 vccd1
+ _14456_/D sky130_fd_sc_hd__o221a_1
XFILLER_203_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _13976_/Q _08095_/A _08190_/X _08097_/A _08184_/X vssd1 vssd1 vccd1 vccd1
+ _13976_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07142_ _14492_/Q _07136_/X _06817_/X _07137_/X _07139_/X vssd1 vssd1 vccd1 vccd1
+ _14492_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07073_ _08259_/A vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__buf_2
XFILLER_192_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput377 _12214_/X vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__clkbuf_2
Xoutput388 _12224_/X vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput399 _12199_/X vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07975_ _08000_/A vssd1 vssd1 vccd1 vccd1 _07975_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09714_ _10077_/B vssd1 vssd1 vccd1 vccd1 _10058_/B sky130_fd_sc_hd__inv_2
X_06926_ _06935_/A _06926_/B vssd1 vssd1 vccd1 vccd1 _14582_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09642_/X _09644_/X _09642_/X _09644_/X vssd1 vssd1 vccd1 vccd1 _09645_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06857_ _06857_/A vssd1 vssd1 vccd1 vccd1 _06857_/X sky130_fd_sc_hd__buf_1
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09576_ _09586_/A _12367_/X vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__and2_2
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06788_ _08945_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08930_/A vssd1 vssd1 vccd1 vccd1 _08527_/X sky130_fd_sc_hd__clkbuf_4
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _13834_/Q _08452_/X _08243_/X _08453_/X _08457_/X vssd1 vssd1 vccd1 vccd1
+ _13834_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07467_/A sky130_fd_sc_hd__inv_2
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08389_ _08389_/A vssd1 vssd1 vccd1 vccd1 _08389_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10420_ _10415_/Y _10242_/X _10416_/Y _10245_/X _10419_/X vssd1 vssd1 vccd1 vccd1
+ _10421_/D sky130_fd_sc_hd__o221a_1
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _13861_/Q vssd1 vssd1 vccd1 vccd1 _10351_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13070_ _13069_/X _12614_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__mux2_1
X_10282_ _14366_/Q vssd1 vssd1 vccd1 vccd1 _10282_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12021_ _12019_/Y _10234_/A _12020_/Y _10237_/A vssd1 vssd1 vccd1 vccd1 _12021_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13972_ _14095_/CLK _13972_/D vssd1 vssd1 vccd1 vccd1 _13972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12923_ _12541_/X _12922_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12854_ _12524_/X _12853_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12854_/X sky130_fd_sc_hd__mux2_1
XPHY_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11805_ _14359_/Q vssd1 vssd1 vccd1 vccd1 _11805_/Y sky130_fd_sc_hd__inv_2
XPHY_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _09528_/X _12784_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__mux2_1
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14524_ _14637_/CLK _14524_/D vssd1 vssd1 vccd1 vccd1 _14524_/Q sky130_fd_sc_hd__dfxtp_1
X_11736_ _14474_/Q vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__inv_2
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14455_ _14470_/CLK _14455_/D vssd1 vssd1 vccd1 vccd1 _14455_/Q sky130_fd_sc_hd__dfxtp_2
X_11667_ _13221_/Q _11485_/X _14044_/Q _11663_/X _11666_/X vssd1 vssd1 vccd1 vccd1
+ _11667_/X sky130_fd_sc_hd__a221o_4
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ _14188_/CLK _13406_/D vssd1 vssd1 vccd1 vccd1 _13406_/Q sky130_fd_sc_hd__dfxtp_1
X_10618_ _10616_/Y _10455_/X _10617_/Y _10458_/X vssd1 vssd1 vccd1 vccd1 _10618_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _14238_/Q _11406_/X _14433_/Q _11407_/X _11597_/X vssd1 vssd1 vccd1 vccd1
+ _11631_/B sky130_fd_sc_hd__a221oi_2
X_14386_ _14495_/CLK _14386_/D vssd1 vssd1 vccd1 vccd1 _14386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ _13584_/Q vssd1 vssd1 vccd1 vccd1 _10549_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13337_ _13368_/CLK _13337_/D vssd1 vssd1 vccd1 vccd1 _13337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13268_ _14639_/CLK _13268_/D vssd1 vssd1 vccd1 vccd1 _13268_/Q sky130_fd_sc_hd__dfxtp_2
X_12219_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13199_ _14071_/CLK _13199_/D vssd1 vssd1 vccd1 vccd1 _13199_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07760_ _07772_/A vssd1 vssd1 vccd1 vccd1 _07760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06711_ _09519_/A vssd1 vssd1 vccd1 vccd1 _09457_/A sky130_fd_sc_hd__buf_4
XFILLER_65_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07691_ _14215_/Q _07687_/X _07392_/X _07688_/X _07684_/X vssd1 vssd1 vccd1 vccd1
+ _14215_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09430_ _09432_/A _12991_/X vssd1 vssd1 vccd1 vccd1 _13310_/D sky130_fd_sc_hd__and2_1
X_06642_ _06636_/X _06641_/X _06636_/X _06641_/X vssd1 vssd1 vccd1 vccd1 _06642_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09364_/A _12831_/X vssd1 vssd1 vccd1 vccd1 _13366_/D sky130_fd_sc_hd__and2_1
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06573_ _06573_/A vssd1 vssd1 vccd1 vccd1 _06573_/X sky130_fd_sc_hd__buf_1
XFILLER_185_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08312_ _13915_/Q _08310_/X _08150_/X _08311_/X _08305_/X vssd1 vssd1 vccd1 vccd1
+ _13915_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09292_ _13413_/Q _09285_/X _08117_/A _09287_/X _09290_/X vssd1 vssd1 vccd1 vccd1
+ _13413_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_12 _11354_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_23 _09457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A vssd1 vssd1 vccd1 vccd1 _08243_/X sky130_fd_sc_hd__buf_4
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_34 _06801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_45 _07476_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_56 _07771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 _08099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08174_ _08174_/A vssd1 vssd1 vccd1 vccd1 _08174_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_78 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_89 _08886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07125_ _14502_/Q _07119_/X _06781_/X _07120_/X _07122_/X vssd1 vssd1 vccd1 vccd1
+ _14502_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07056_ _14538_/Q _07052_/X _06793_/X _07053_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _14538_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07958_ _14091_/Q _07955_/X _07809_/X _07957_/X _07946_/X vssd1 vssd1 vccd1 vccd1
+ _14091_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06909_ _14586_/Q vssd1 vssd1 vccd1 vccd1 _06909_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07889_ _14127_/Q _07882_/X _07712_/X _07884_/X _07886_/X vssd1 vssd1 vccd1 vccd1
+ _14127_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09628_ _09622_/X _09627_/X _09622_/X _09627_/X vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ _09557_/X _09556_/X _13271_/Q _09558_/X vssd1 vssd1 vccd1 vccd1 _13239_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _13296_/Q _12569_/X input39/X vssd1 vssd1 vccd1 vccd1 _12570_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11521_ _13846_/Q vssd1 vssd1 vccd1 vccd1 _11521_/Y sky130_fd_sc_hd__inv_2
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14240_ _14633_/CLK _14240_/D vssd1 vssd1 vccd1 vccd1 _14240_/Q sky130_fd_sc_hd__dfxtp_1
X_11452_ _11448_/Y _11449_/X _11450_/Y _11451_/X vssd1 vssd1 vccd1 vccd1 _11452_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ _14486_/Q vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ _14173_/CLK _14171_/D vssd1 vssd1 vccd1 vccd1 _14171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11383_ _13602_/Q vssd1 vssd1 vccd1 vccd1 _11383_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10334_ _14133_/Q vssd1 vssd1 vccd1 vccd1 _10334_/Y sky130_fd_sc_hd__inv_2
X_13122_ _13121_/X _12639_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13053_ _12606_/X _13052_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10265_ _13742_/Q vssd1 vssd1 vccd1 vccd1 _10265_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12004_ _12002_/Y _10188_/A _12003_/Y _10191_/A vssd1 vssd1 vccd1 vccd1 _12004_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10196_ _13500_/Q vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13955_ _13996_/CLK _13955_/D vssd1 vssd1 vccd1 vccd1 _13955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12906_ _12537_/X _12905_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12906_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13886_ _14100_/CLK _13886_/D vssd1 vssd1 vccd1 vccd1 _13886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12837_ _12520_/X _12836_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12837_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12768_ _09519_/X input353/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12768_/X sky130_fd_sc_hd__mux2_1
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14507_ _14627_/CLK _14507_/D vssd1 vssd1 vccd1 vccd1 _14507_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _13570_/Q _11664_/X _13811_/Q _11665_/X vssd1 vssd1 vccd1 vccd1 _11719_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12699_ _09597_/X _12698_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13191_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14438_ _14481_/CLK _14438_/D vssd1 vssd1 vccd1 vccd1 _14438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput21 io_in[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xinput32 io_in[3] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_1
XFILLER_15_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput43 la_data_in[103] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
XFILLER_174_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput54 la_data_in[113] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_1
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14369_ _14633_/CLK _14369_/D vssd1 vssd1 vccd1 vccd1 _14369_/Q sky130_fd_sc_hd__dfxtp_1
Xinput65 la_data_in[123] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_1
Xinput76 la_data_in[18] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
XFILLER_7_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput87 la_data_in[28] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_1
XFILLER_171_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput98 la_data_in[38] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_2
XFILLER_118_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _08930_/A vssd1 vssd1 vccd1 vccd1 _08930_/X sky130_fd_sc_hd__buf_6
XFILLER_63_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08861_ _08869_/A vssd1 vssd1 vccd1 vccd1 _08861_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07812_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07812_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater611 _12505_/S vssd1 vssd1 vccd1 vccd1 _12502_/S sky130_fd_sc_hd__buf_8
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08792_ _08792_/A vssd1 vssd1 vccd1 vccd1 _08792_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater622 _12368_/S vssd1 vssd1 vccd1 vccd1 _12407_/S sky130_fd_sc_hd__buf_6
XFILLER_211_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater633 _12888_/S vssd1 vssd1 vccd1 vccd1 _13144_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater644 _14495_/CLK vssd1 vssd1 vccd1 vccd1 _14627_/CLK sky130_fd_sc_hd__buf_12
XFILLER_6_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater655 _14178_/CLK vssd1 vssd1 vccd1 vccd1 _14529_/CLK sky130_fd_sc_hd__buf_12
X_07743_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07743_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater666 _14047_/CLK vssd1 vssd1 vccd1 vccd1 _14121_/CLK sky130_fd_sc_hd__buf_6
XFILLER_113_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater677 _13996_/CLK vssd1 vssd1 vccd1 vccd1 _13877_/CLK sky130_fd_sc_hd__buf_12
XPHY_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater688 _12655_/S vssd1 vssd1 vccd1 vccd1 _12659_/S sky130_fd_sc_hd__buf_8
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater699 _13141_/S vssd1 vssd1 vccd1 vccd1 _13133_/S sky130_fd_sc_hd__buf_8
X_07674_ _09336_/A vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06625_ _06626_/A vssd1 vssd1 vccd1 vccd1 _06625_/Y sky130_fd_sc_hd__inv_2
X_09413_ _09413_/A _13067_/X vssd1 vssd1 vccd1 vccd1 _13323_/D sky130_fd_sc_hd__and2_1
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09344_ _09345_/A _12907_/X vssd1 vssd1 vccd1 vccd1 _13379_/D sky130_fd_sc_hd__and2_1
X_06556_ _06558_/A vssd1 vssd1 vccd1 vccd1 _06556_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09275_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ _13962_/Q _08221_/X _08128_/X _08222_/X _08223_/X vssd1 vssd1 vccd1 vccd1
+ _13962_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _13990_/Q _08149_/X _07852_/X _08151_/X _08147_/X vssd1 vssd1 vccd1 vccd1
+ _13990_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07108_ _14513_/Q _07102_/X _07031_/X _07104_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _14513_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08088_ _14015_/Q _08025_/A _07800_/X _08027_/A _08083_/X vssd1 vssd1 vccd1 vccd1
+ _14015_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07039_ _14549_/Q _07035_/X _06753_/X _07036_/X _07038_/X vssd1 vssd1 vccd1 vccd1
+ _14549_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _13353_/Q _09967_/B _13353_/Q _09967_/B vssd1 vssd1 vccd1 vccd1 _10050_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_7413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _14169_/CLK _13740_/D vssd1 vssd1 vccd1 vccd1 _13740_/Q sky130_fd_sc_hd__dfxtp_1
X_10952_ _11424_/A vssd1 vssd1 vccd1 vccd1 _10952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13671_ _14071_/CLK _13671_/D vssd1 vssd1 vccd1 vccd1 _13671_/Q sky130_fd_sc_hd__dfxtp_1
X_10883_ _13670_/Q vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ _09844_/Y _13333_/Q _12650_/S vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__mux2_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _13289_/Q _12552_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11504_ _11502_/Y _11459_/X _11503_/Y _11461_/X vssd1 vssd1 vccd1 vccd1 _11504_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _12483_/X _06964_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__mux2_2
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14305_/CLK _14223_/D vssd1 vssd1 vccd1 vccd1 _14223_/Q sky130_fd_sc_hd__dfxtp_1
X_11435_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11366_ _11364_/Y _11178_/X _11365_/Y _11180_/X vssd1 vssd1 vccd1 vccd1 _11366_/X
+ sky130_fd_sc_hd__o22a_1
X_14154_ _14305_/CLK _14154_/D vssd1 vssd1 vccd1 vccd1 _14154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10317_ _10315_/Y _10195_/X _10316_/Y _10198_/X vssd1 vssd1 vccd1 vccd1 _10317_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _12631_/X _13104_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14085_ _14178_/CLK _14085_/D vssd1 vssd1 vccd1 vccd1 _14085_/Q sky130_fd_sc_hd__dfxtp_1
X_11297_ _14387_/Q vssd1 vssd1 vccd1 vccd1 _11297_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10248_ _10248_/A vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__clkbuf_2
X_13036_ _12598_/X input349/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10179_ _13741_/Q vssd1 vssd1 vccd1 vccd1 _10179_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _14095_/CLK _13938_/D vssd1 vssd1 vccd1 vccd1 _13938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13869_ _14107_/CLK _13869_/D vssd1 vssd1 vccd1 vccd1 _13869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07390_ _14373_/Q _07387_/X _07388_/X _07389_/X _07385_/X vssd1 vssd1 vccd1 vccd1
+ _14373_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09060_ _09060_/A vssd1 vssd1 vccd1 vccd1 _09060_/X sky130_fd_sc_hd__buf_4
XFILLER_31_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08011_ _08017_/A vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09962_ _09886_/A _09886_/B _09961_/Y vssd1 vssd1 vccd1 vccd1 _09962_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08913_ _13608_/Q _08905_/X _08912_/X _08907_/X _08910_/X vssd1 vssd1 vccd1 vccd1
+ _13608_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09893_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__or2_1
XFILLER_115_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08868_/A vssd1 vssd1 vccd1 vccd1 _08844_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _08792_/A vssd1 vssd1 vccd1 vccd1 _08775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07726_ _08117_/A vssd1 vssd1 vccd1 vccd1 _07726_/X sky130_fd_sc_hd__buf_4
XPHY_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07657_ _14235_/Q _07653_/X _07341_/X _07654_/X _07650_/X vssd1 vssd1 vccd1 vccd1
+ _14235_/D sky130_fd_sc_hd__o221a_1
XFILLER_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06608_ _06608_/A vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__clkbuf_4
X_07588_ _14272_/Q _07580_/X _07345_/X _07581_/X _07585_/X vssd1 vssd1 vccd1 vccd1
+ _14272_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09327_ _09327_/A vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06539_ _06541_/A vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__buf_4
XFILLER_179_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08209_ _13970_/Q _08198_/X _08105_/X _08201_/X _08204_/X vssd1 vssd1 vccd1 vccd1
+ _13970_/D sky130_fd_sc_hd__o221a_1
X_09189_ _09189_/A vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11220_ _14151_/Q vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11151_ _11146_/Y _10973_/X _11147_/Y _10975_/X _11150_/X vssd1 vssd1 vccd1 vccd1
+ _11158_/C sky130_fd_sc_hd__o221a_1
XFILLER_46_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ _10107_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__or2_1
XFILLER_81_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11082_ _11080_/Y _10927_/X _11081_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _11082_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput200 la_oenb[14] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__buf_1
XPHY_7221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput211 la_oenb[24] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_1
XFILLER_42_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _13370_/Q _09998_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _10033_/X sky130_fd_sc_hd__o21a_1
Xinput222 la_oenb[34] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_1
XFILLER_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput233 la_oenb[44] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_1
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 la_oenb[54] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_1
XPHY_7265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput255 la_oenb[64] vssd1 vssd1 vccd1 vccd1 _12283_/S sky130_fd_sc_hd__buf_1
XPHY_7276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput266 la_oenb[74] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_hd__buf_1
XPHY_7287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput277 la_oenb[84] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_hd__buf_1
XPHY_7298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput288 la_oenb[94] vssd1 vssd1 vccd1 vccd1 input288/X sky130_fd_sc_hd__buf_1
XFILLER_64_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput299 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _06503_/C sky130_fd_sc_hd__clkbuf_1
XPHY_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ _13498_/Q vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13723_ _14183_/CLK _13723_/D vssd1 vssd1 vccd1 vccd1 _13723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10935_ _11407_/A vssd1 vssd1 vccd1 vccd1 _10935_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ _14056_/CLK _13654_/D vssd1 vssd1 vccd1 vccd1 _13654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ _10861_/Y _10725_/X _10862_/Y _10727_/X _10865_/X vssd1 vssd1 vccd1 vccd1
+ _10879_/B sky130_fd_sc_hd__o221a_4
XFILLER_182_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _09856_/Y _13326_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12605_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _14178_/CLK _13585_/D vssd1 vssd1 vccd1 vccd1 _13585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _10797_/A _10797_/B _10797_/C _10797_/D vssd1 vssd1 vccd1 vccd1 _10797_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12536_ _13380_/Q _10024_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12536_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12467_ _12509_/X _06943_/X _12467_/S vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _14325_/CLK _14206_/D vssd1 vssd1 vccd1 vccd1 _14206_/Q sky130_fd_sc_hd__dfxtp_1
X_11418_ _13844_/Q vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12398_ _13221_/Q _06611_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12398_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14137_ _14139_/CLK _14137_/D vssd1 vssd1 vccd1 vccd1 _14137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11349_ _13484_/Q vssd1 vssd1 vccd1 vccd1 _11349_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14068_ _14071_/CLK _14068_/D vssd1 vssd1 vccd1 vccd1 _14068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13019_ _12588_/X _13018_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13019_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06890_ _06880_/X _12291_/X _06889_/Y _06883_/X vssd1 vssd1 vccd1 vccd1 _06891_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08560_ _08965_/A vssd1 vssd1 vccd1 vccd1 _08560_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07511_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07511_/X sky130_fd_sc_hd__clkbuf_2
X_08491_ _13817_/Q _08486_/X _08490_/X _08488_/X _08480_/X vssd1 vssd1 vccd1 vccd1
+ _13817_/D sky130_fd_sc_hd__o221a_1
XFILLER_169_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ _09336_/A vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09112_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ _13550_/Q _09039_/X _08962_/X _09040_/X _09036_/X vssd1 vssd1 vccd1 vccd1
+ _13550_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _13296_/Q _09943_/Y _09891_/B vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09876_ _13292_/Q vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__inv_2
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08827_ _08827_/A vssd1 vssd1 vccd1 vccd1 _08827_/X sky130_fd_sc_hd__buf_4
XPHY_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08792_/A vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07709_ _14207_/Q _07704_/X _07708_/X _07706_/X _07698_/X vssd1 vssd1 vccd1 vccd1
+ _14207_/D sky130_fd_sc_hd__o221a_1
XPHY_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08689_ _08723_/A vssd1 vssd1 vccd1 vccd1 _08689_/X sky130_fd_sc_hd__buf_2
XPHY_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10720_ _11430_/A vssd1 vssd1 vccd1 vccd1 _10720_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10651_ _13392_/Q _10568_/X _13704_/Q _10440_/X vssd1 vssd1 vccd1 vccd1 _10651_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10582_ _13546_/Q _10471_/X _13787_/Q _10473_/X vssd1 vssd1 vccd1 vccd1 _10582_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13370_ _13370_/CLK _13370_/D vssd1 vssd1 vccd1 vccd1 _13370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ _10298_/Y _14522_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12321_/X sky130_fd_sc_hd__mux2_4
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12252_ _12033_/Y _13353_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _11439_/A vssd1 vssd1 vccd1 vccd1 _11203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12183_ vssd1 vssd1 vccd1 vccd1 _12183_/HI _12183_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11134_ _13994_/Q vssd1 vssd1 vccd1 vccd1 _11134_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11065_ _13595_/Q vssd1 vssd1 vccd1 vccd1 _11065_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10016_ _10016_/A vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__inv_2
XFILLER_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11957_/Y _10178_/A _11960_/X _11963_/X _11966_/X vssd1 vssd1 vccd1 vccd1
+ _11989_/C sky130_fd_sc_hd__o2111a_4
XPHY_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13706_ _14183_/CLK _13706_/D vssd1 vssd1 vccd1 vccd1 _13706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ _10916_/Y _10749_/X _10917_/Y _10751_/X vssd1 vssd1 vccd1 vccd1 _10918_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _11896_/Y _10234_/A _11897_/Y _10237_/A vssd1 vssd1 vccd1 vccd1 _11898_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ _14071_/CLK _13637_/D vssd1 vssd1 vccd1 vccd1 _13637_/Q sky130_fd_sc_hd__dfxtp_1
X_10849_ _13754_/Q vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13568_ _14121_/CLK _13568_/D vssd1 vssd1 vccd1 vccd1 _13568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12519_ _13365_/Q _10044_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12519_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13499_ _14173_/CLK _13499_/D vssd1 vssd1 vccd1 vccd1 _13499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput504 _12135_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput515 _12145_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput526 _12155_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput537 _12165_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__clkbuf_2
Xoutput548 _12175_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__clkbuf_2
Xoutput559 _12185_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07991_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09730_ _06869_/A _09729_/X _06869_/A _09729_/X vssd1 vssd1 vccd1 vccd1 _09730_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06942_ _14577_/Q vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__inv_2
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _06869_/X _09660_/Y _06869_/X _09660_/Y vssd1 vssd1 vccd1 vccd1 _09661_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06873_ _06857_/X _12287_/X _06872_/Y _06861_/X vssd1 vssd1 vccd1 vccd1 _06874_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08612_ _08637_/A vssd1 vssd1 vccd1 vccd1 _08612_/X sky130_fd_sc_hd__buf_1
XFILLER_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09592_ _09583_/X _09591_/X _13258_/Q _09584_/X vssd1 vssd1 vccd1 vccd1 _13226_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08543_ _13798_/Q _08540_/X _08541_/X _08542_/X _08538_/X vssd1 vssd1 vccd1 vccd1
+ _13798_/D sky130_fd_sc_hd__o221a_1
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08474_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07356_ _08144_/A vssd1 vssd1 vccd1 vccd1 _07356_/X sky130_fd_sc_hd__buf_2
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07287_ _07301_/A vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09026_ _13560_/Q _09022_/X _08935_/X _09023_/X _09019_/X vssd1 vssd1 vccd1 vccd1
+ _13560_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09928_ _09926_/A _09926_/B _09927_/Y vssd1 vssd1 vccd1 vccd1 _09928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09859_ _13309_/Q vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__inv_2
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12528_/X _12869_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12870_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_102 _09383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11816_/Y _11689_/X _11817_/Y _11691_/X _11820_/X vssd1 vssd1 vccd1 vccd1
+ _11822_/D sky130_fd_sc_hd__o221a_1
XPHY_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_113 _11457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _11139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _11293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_146 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_157 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14621_/CLK _14540_/D vssd1 vssd1 vccd1 vccd1 _14540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11752_ _13890_/Q vssd1 vssd1 vccd1 vccd1 _11752_/Y sky130_fd_sc_hd__inv_2
XPHY_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 input333/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10703_ _13751_/Q vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__inv_2
XPHY_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14471_ _14611_/CLK _14471_/D vssd1 vssd1 vccd1 vccd1 _14471_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11683_ _11683_/A vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__buf_2
XPHY_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13422_ _14056_/CLK _13422_/D vssd1 vssd1 vccd1 vccd1 _13422_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10634_ _14256_/Q vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13353_ _14639_/CLK _13353_/D vssd1 vssd1 vccd1 vccd1 _13353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10565_ _13624_/Q vssd1 vssd1 vccd1 vccd1 _10565_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12304_ _11118_/Y _14539_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12304_/X sky130_fd_sc_hd__mux2_2
X_13284_ _14538_/CLK _13284_/D vssd1 vssd1 vccd1 vccd1 _13284_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10496_ _14175_/Q vssd1 vssd1 vccd1 vccd1 _10496_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ _12235_/A vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12166_ vssd1 vssd1 vccd1 vccd1 _12166_/HI _12166_/LO sky130_fd_sc_hd__conb_1
XFILLER_116_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11117_ _11098_/X _11117_/B _11117_/C _11117_/D vssd1 vssd1 vccd1 vccd1 _11118_/D
+ sky130_fd_sc_hd__and4b_1
X_12097_ vssd1 vssd1 vccd1 vccd1 _12097_/HI _12097_/LO sky130_fd_sc_hd__conb_1
XFILLER_211_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11048_ _11046_/Y _10942_/X _11047_/Y _10944_/X vssd1 vssd1 vccd1 vccd1 _11048_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12999_ _12578_/X _12998_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08190_ _08190_/A vssd1 vssd1 vccd1 vccd1 _08190_/X sky130_fd_sc_hd__buf_4
XFILLER_203_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ _14493_/Q _07136_/X _06814_/X _07137_/X _07139_/X vssd1 vssd1 vccd1 vccd1
+ _14493_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07072_ _14529_/Q _07069_/X _06825_/X _07070_/X _07071_/X vssd1 vssd1 vccd1 vccd1
+ _14529_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput378 _12215_/X vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput389 _12225_/X vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07974_ _07999_/A vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09713_ _10128_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__or2_1
XFILLER_45_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06925_ _06919_/X _12300_/X _06924_/Y _06921_/X vssd1 vssd1 vccd1 vccd1 _06926_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09644_ _14566_/Q _09643_/X _14566_/Q _09643_/X vssd1 vssd1 vccd1 vccd1 _09644_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06856_ _09650_/A vssd1 vssd1 vccd1 vccd1 _06857_/A sky130_fd_sc_hd__buf_1
XFILLER_167_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09575_ _09588_/A vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__buf_1
XFILLER_43_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06787_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06787_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08526_ _08552_/A vssd1 vssd1 vccd1 vccd1 _08526_/X sky130_fd_sc_hd__clkbuf_2
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08457_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07408_ _07558_/A _11671_/A vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__or2_2
XFILLER_127_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08388_ _08388_/A vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07339_ _08126_/A vssd1 vssd1 vccd1 vccd1 _07339_/X sky130_fd_sc_hd__buf_2
XFILLER_32_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _13744_/Q vssd1 vssd1 vccd1 vccd1 _10350_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ _09009_/A vssd1 vssd1 vccd1 vccd1 _09009_/X sky130_fd_sc_hd__buf_4
XFILLER_178_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10281_ _14600_/Q vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ _14286_/Q vssd1 vssd1 vccd1 vccd1 _12020_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13971_ _14095_/CLK _13971_/D vssd1 vssd1 vccd1 vccd1 _13971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12922_ _12541_/X _12921_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12853_ _12524_/X _12852_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11804_ _14515_/Q vssd1 vssd1 vccd1 vccd1 _11804_/Y sky130_fd_sc_hd__inv_2
XPHY_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12784_ _09528_/X input348/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__mux2_1
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14523_ _14637_/CLK _14523_/D vssd1 vssd1 vccd1 vccd1 _14523_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11735_ _13492_/Q vssd1 vssd1 vccd1 vccd1 _11735_/Y sky130_fd_sc_hd__inv_2
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _14470_/CLK _14454_/D vssd1 vssd1 vccd1 vccd1 _14454_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _13569_/Q _11664_/X _13810_/Q _11665_/X vssd1 vssd1 vccd1 vccd1 _11666_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _14188_/CLK _13405_/D vssd1 vssd1 vccd1 vccd1 _13405_/Q sky130_fd_sc_hd__dfxtp_1
X_10617_ _14100_/Q vssd1 vssd1 vccd1 vccd1 _10617_/Y sky130_fd_sc_hd__inv_2
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14385_ _14495_/CLK _14385_/D vssd1 vssd1 vccd1 vccd1 _14385_/Q sky130_fd_sc_hd__dfxtp_1
X_11597_ _13412_/Q _11514_/X _13724_/Q _11408_/X vssd1 vssd1 vccd1 vccd1 _11597_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ _13352_/CLK _13336_/D vssd1 vssd1 vccd1 vccd1 _13336_/Q sky130_fd_sc_hd__dfxtp_1
X_10548_ _14293_/Q vssd1 vssd1 vccd1 vccd1 _10548_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13267_ _14639_/CLK _13267_/D vssd1 vssd1 vccd1 vccd1 _13267_/Q sky130_fd_sc_hd__dfxtp_2
X_10479_ _14331_/Q vssd1 vssd1 vccd1 vccd1 _10479_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12218_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13198_ _13352_/CLK _13198_/D vssd1 vssd1 vccd1 vccd1 _13198_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12149_ vssd1 vssd1 vccd1 vccd1 _12149_/HI _12149_/LO sky130_fd_sc_hd__conb_1
XFILLER_155_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06710_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__buf_2
XFILLER_42_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07690_ _14216_/Q _07687_/X _07471_/X _07688_/X _07684_/X vssd1 vssd1 vccd1 vccd1
+ _14216_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06641_ _06637_/Y _06640_/X _06637_/Y _06640_/X vssd1 vssd1 vccd1 vccd1 _06641_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09360_ _09364_/A _12891_/X vssd1 vssd1 vccd1 vccd1 _13367_/D sky130_fd_sc_hd__and2_1
X_06572_ _06611_/A vssd1 vssd1 vccd1 vccd1 _06573_/A sky130_fd_sc_hd__inv_2
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08311_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09291_ _13414_/Q _09285_/X _09009_/X _09287_/X _09290_/X vssd1 vssd1 vccd1 vccd1
+ _13414_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_13 _11465_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08242_ _13952_/Q _08237_/X _08155_/X _08238_/X _08239_/X vssd1 vssd1 vccd1 vccd1
+ _13952_/D sky130_fd_sc_hd__o221a_1
XANTENNA_24 _08217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_35 _08181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_46 _07532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_57 _07771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 _08099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _13984_/Q _08161_/X _08171_/X _08163_/X _08172_/X vssd1 vssd1 vccd1 vccd1
+ _13984_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_79 _08181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07124_ _14503_/Q _07119_/X _06778_/X _07120_/X _07122_/X vssd1 vssd1 vccd1 vccd1
+ _14503_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07055_ _14539_/Q _07052_/X _06789_/X _07053_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _14539_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ _07957_/A vssd1 vssd1 vccd1 vccd1 _07957_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06908_ _06917_/A _06908_/B vssd1 vssd1 vccd1 vccd1 _14587_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07888_ _14128_/Q _07882_/X _07710_/X _07884_/X _07886_/X vssd1 vssd1 vccd1 vccd1
+ _14128_/D sky130_fd_sc_hd__o221a_1
XFILLER_186_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09627_ _09623_/X _09626_/X _09623_/X _09626_/X vssd1 vssd1 vccd1 vccd1 _09627_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06839_ _14603_/Q _06823_/X _06837_/X _06532_/A _06838_/X vssd1 vssd1 vccd1 vccd1
+ _14603_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09558_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09558_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08509_ _13810_/Q _08500_/X _08508_/X _08503_/X _08497_/X vssd1 vssd1 vccd1 vccd1
+ _13810_/D sky130_fd_sc_hd__o221a_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ _13270_/Q _09486_/X _12265_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _13270_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11520_ _11518_/Y _11414_/X _11519_/Y _11416_/X vssd1 vssd1 vccd1 vccd1 _11520_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11451_ _11451_/A vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _13195_/Q _10276_/X _14018_/Q _10203_/X _10401_/X vssd1 vssd1 vccd1 vccd1
+ _10402_/X sky130_fd_sc_hd__a221o_2
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14170_ _14325_/CLK _14170_/D vssd1 vssd1 vccd1 vccd1 _14170_/Q sky130_fd_sc_hd__dfxtp_1
X_11382_ _14311_/Q vssd1 vssd1 vccd1 vccd1 _11382_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13121_ _12639_/X _13120_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ _13899_/Q vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _12606_/X input359/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10264_ _13937_/Q vssd1 vssd1 vccd1 vccd1 _10264_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12003_ _14130_/Q vssd1 vssd1 vccd1 vccd1 _12003_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10195_ _10195_/A vssd1 vssd1 vccd1 vccd1 _10195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13954_ _14107_/CLK _13954_/D vssd1 vssd1 vccd1 vccd1 _13954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12905_ _12537_/X _12904_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13885_ _14100_/CLK _13885_/D vssd1 vssd1 vccd1 vccd1 _13885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12836_ _12520_/X input334/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12767_ _09509_/X _12766_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13222_/D sky130_fd_sc_hd__mux2_1
XFILLER_206_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14506_ _14627_/CLK _14506_/D vssd1 vssd1 vccd1 vccd1 _14506_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _11708_/Y _11646_/X _11711_/X _11714_/X _11717_/X vssd1 vssd1 vccd1 vccd1
+ _11740_/C sky130_fd_sc_hd__o2111a_4
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12698_ _09597_/X _12697_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12698_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14437_ _14527_/CLK _14437_/D vssd1 vssd1 vccd1 vccd1 _14437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
X_11649_ _13888_/Q vssd1 vssd1 vccd1 vccd1 _11649_/Y sky130_fd_sc_hd__inv_2
Xinput22 io_in[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 io_in[4] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
Xinput44 la_data_in[104] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
XFILLER_176_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14368_ _14633_/CLK _14368_/D vssd1 vssd1 vccd1 vccd1 _14368_/Q sky130_fd_sc_hd__dfxtp_1
Xinput55 la_data_in[114] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
XFILLER_102_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput66 la_data_in[124] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_1
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput77 la_data_in[19] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_1
XFILLER_85_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput88 la_data_in[29] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_1
X_13319_ _14114_/CLK _13319_/D vssd1 vssd1 vccd1 vccd1 _13319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput99 la_data_in[39] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_2
XFILLER_171_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14299_ _14305_/CLK _14299_/D vssd1 vssd1 vccd1 vccd1 _14299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ _08868_/A vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07811_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07811_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater612 _12603_/S vssd1 vssd1 vccd1 vccd1 _12601_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08791_ _13670_/Q _08783_/X _08549_/X _08784_/X _08786_/X vssd1 vssd1 vccd1 vccd1
+ _13670_/D sky130_fd_sc_hd__o221a_1
Xrepeater623 _09601_/X vssd1 vssd1 vccd1 vccd1 _12368_/S sky130_fd_sc_hd__buf_8
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater634 _09796_/X vssd1 vssd1 vccd1 vccd1 _13176_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_211_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater645 _14611_/CLK vssd1 vssd1 vccd1 vccd1 _14495_/CLK sky130_fd_sc_hd__buf_8
XFILLER_22_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater656 _14139_/CLK vssd1 vssd1 vccd1 vccd1 _14178_/CLK sky130_fd_sc_hd__buf_12
X_07742_ _08132_/A vssd1 vssd1 vccd1 vccd1 _07742_/X sky130_fd_sc_hd__buf_4
Xrepeater667 _14119_/CLK vssd1 vssd1 vccd1 vccd1 _14047_/CLK sky130_fd_sc_hd__buf_12
XFILLER_6_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater678 _14114_/CLK vssd1 vssd1 vccd1 vccd1 _13996_/CLK sky130_fd_sc_hd__buf_12
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater689 _12645_/S vssd1 vssd1 vccd1 vccd1 _12655_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07673_ _14225_/Q _07669_/X _07367_/X _07670_/X _07666_/X vssd1 vssd1 vccd1 vccd1
+ _14225_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09412_ _09413_/A _13063_/X vssd1 vssd1 vccd1 vccd1 _13324_/D sky130_fd_sc_hd__and2_1
XFILLER_168_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06624_ _06699_/A _06623_/X _06699_/A _06623_/X vssd1 vssd1 vccd1 vccd1 _06624_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09343_ _09345_/A _12903_/X vssd1 vssd1 vccd1 vccd1 _13380_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06555_ _08917_/A _08940_/A _06553_/Y _06554_/Y vssd1 vssd1 vccd1 vccd1 _06562_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _09326_/A vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _13963_/Q _08221_/X _08126_/X _08222_/X _08223_/X vssd1 vssd1 vccd1 vccd1
+ _13963_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08156_ _13991_/Q _08149_/X _08155_/X _08151_/X _08147_/X vssd1 vssd1 vccd1 vccd1
+ _13991_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07107_ _14514_/Q _07102_/X _06738_/X _07104_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _14514_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08087_ _14016_/Q _08025_/A _07798_/X _08027_/A _08083_/X vssd1 vssd1 vccd1 vccd1
+ _14016_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07038_ _07071_/A vssd1 vssd1 vccd1 vccd1 _07038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _08989_/A _08989_/B _08989_/C _08989_/D vssd1 vssd1 vccd1 vccd1 _10204_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_25_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _13990_/Q vssd1 vssd1 vccd1 vccd1 _10951_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13670_ _14071_/CLK _13670_/D vssd1 vssd1 vccd1 vccd1 _13670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10882_ _13436_/Q vssd1 vssd1 vccd1 vccd1 _10882_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _13334_/Q _12620_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__mux2_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _09957_/Y _13289_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12552_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _14469_/Q vssd1 vssd1 vccd1 vccd1 _11503_/Y sky130_fd_sc_hd__inv_2
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12483_ _12482_/X _06964_/Y _12486_/S vssd1 vssd1 vccd1 vccd1 _12483_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14222_ _14470_/CLK _14222_/D vssd1 vssd1 vccd1 vccd1 _14222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11434_ _14507_/Q vssd1 vssd1 vccd1 vccd1 _11434_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14153_ _14595_/CLK _14153_/D vssd1 vssd1 vccd1 vccd1 _14153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11365_ _13882_/Q vssd1 vssd1 vccd1 vccd1 _11365_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _12631_/X input331/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13104_/X sky130_fd_sc_hd__mux2_1
X_10316_ _13502_/Q vssd1 vssd1 vccd1 vccd1 _10316_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14084_ _14291_/CLK _14084_/D vssd1 vssd1 vccd1 vccd1 _14084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11296_ _14621_/Q vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13035_ _12596_/X _13034_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ _11693_/A vssd1 vssd1 vccd1 vccd1 _10248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _10178_/A vssd1 vssd1 vccd1 vccd1 _10178_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13937_ _14095_/CLK _13937_/D vssd1 vssd1 vccd1 vccd1 _13937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13868_ _14107_/CLK _13868_/D vssd1 vssd1 vccd1 vccd1 _13868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12819_ _12516_/X _12818_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12819_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13799_ _14114_/CLK _13799_/D vssd1 vssd1 vccd1 vccd1 _13799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08010_ _14060_/Q _08007_/X _07867_/X _08008_/X _08003_/X vssd1 vssd1 vccd1 vccd1
+ _14060_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _09961_/A vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08912_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__buf_4
XFILLER_8_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09892_ _09892_/A _09946_/A vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__or2_1
XFILLER_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ _13646_/Q _08832_/X _08510_/X _08835_/X _08839_/X vssd1 vssd1 vccd1 vccd1
+ _13646_/D sky130_fd_sc_hd__o221a_1
XFILLER_189_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _13680_/Q _08767_/X _08523_/X _08768_/X _08769_/X vssd1 vssd1 vccd1 vccd1
+ _13680_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07725_ _14201_/Q _07718_/X _07428_/X _07721_/X _07715_/X vssd1 vssd1 vccd1 vccd1
+ _14201_/D sky130_fd_sc_hd__o221a_1
XPHY_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07656_ _14236_/Q _07653_/X _07339_/X _07654_/X _07650_/X vssd1 vssd1 vccd1 vccd1
+ _14236_/D sky130_fd_sc_hd__o221a_1
XPHY_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ _06587_/X _06606_/Y _06587_/X _06606_/Y vssd1 vssd1 vccd1 vccd1 _06608_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07587_ _14273_/Q _07580_/X _07343_/X _07581_/X _07585_/X vssd1 vssd1 vccd1 vccd1
+ _14273_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _09326_/A vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06538_ _06540_/A vssd1 vssd1 vccd1 vccd1 _06538_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09257_ _09257_/A vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08208_ _13971_/Q _08198_/X _08103_/X _08201_/X _08204_/X vssd1 vssd1 vccd1 vccd1
+ _13971_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ _09188_/A vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08139_ _13998_/Q _08136_/X _08137_/X _08138_/X _08134_/X vssd1 vssd1 vccd1 vccd1
+ _13998_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11150_ _11148_/Y _10977_/X _11149_/Y _10979_/X vssd1 vssd1 vccd1 vccd1 _11150_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10101_ _10114_/A _12475_/X vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__nor2_8
XFILLER_27_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11081_ _13635_/Q vssd1 vssd1 vccd1 vccd1 _11081_/Y sky130_fd_sc_hd__inv_2
XPHY_7200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput201 la_oenb[15] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__buf_1
XPHY_7222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _13369_/Q _09996_/B _09997_/A vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__o21a_1
Xinput212 la_oenb[25] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__buf_1
XFILLER_103_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput223 la_oenb[35] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_1
XPHY_7244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 la_oenb[45] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_1
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 la_oenb[55] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_1
XPHY_7266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput256 la_oenb[65] vssd1 vssd1 vccd1 vccd1 _12282_/S sky130_fd_sc_hd__buf_1
XPHY_7277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput267 la_oenb[75] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__buf_1
XPHY_7288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput278 la_oenb[85] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_hd__buf_1
XPHY_7299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput289 la_oenb[95] vssd1 vssd1 vccd1 vccd1 input289/X sky130_fd_sc_hd__buf_1
XFILLER_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11983_ _14168_/Q vssd1 vssd1 vccd1 vccd1 _11983_/Y sky130_fd_sc_hd__inv_2
XPHY_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13722_ _14183_/CLK _13722_/D vssd1 vssd1 vccd1 vccd1 _13722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ _11831_/A vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__buf_4
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13653_ _14056_/CLK _13653_/D vssd1 vssd1 vccd1 vccd1 _13653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10865_ _10863_/Y _10729_/X _10864_/Y _10731_/X vssd1 vssd1 vccd1 vccd1 _10865_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _13311_/Q _12603_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12604_/X sky130_fd_sc_hd__mux2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13584_ _14178_/CLK _13584_/D vssd1 vssd1 vccd1 vccd1 _13584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10777_/X _10796_/B _10796_/C _10796_/D vssd1 vssd1 vccd1 vccd1 _10797_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12535_ _13381_/Q _10027_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12535_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12466_ _12465_/X _06938_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12466_/X sky130_fd_sc_hd__mux2_2
XFILLER_138_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14205_ _14325_/CLK _14205_/D vssd1 vssd1 vccd1 vccd1 _14205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _11413_/Y _11414_/X _11415_/Y _11416_/X vssd1 vssd1 vccd1 vccd1 _11417_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12397_ _12396_/X _13222_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12397_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14136_ _14139_/CLK _14136_/D vssd1 vssd1 vccd1 vccd1 _14136_/Q sky130_fd_sc_hd__dfxtp_1
X_11348_ _14154_/Q vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14067_ _14071_/CLK _14067_/D vssd1 vssd1 vccd1 vccd1 _14067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11279_ _13405_/Q _11278_/X _13717_/Q _11172_/X vssd1 vssd1 vccd1 vccd1 _11279_/X
+ sky130_fd_sc_hd__a22o_2
X_13018_ _13017_/X _12588_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _13018_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07510_ _14315_/Q _07508_/X _07336_/X _07509_/X _07503_/X vssd1 vssd1 vccd1 vccd1
+ _14315_/D sky130_fd_sc_hd__o221a_1
X_08490_ _08822_/A vssd1 vssd1 vccd1 vccd1 _08490_/X sky130_fd_sc_hd__buf_2
XFILLER_93_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07372_ _14379_/Q _07361_/X _07370_/X _07363_/X _07371_/X vssd1 vssd1 vccd1 vccd1
+ _14379_/D sky130_fd_sc_hd__o221a_1
XFILLER_182_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09042_ _13551_/Q _09039_/X _08960_/X _09040_/X _09036_/X vssd1 vssd1 vccd1 vccd1
+ _13551_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09944_ _09889_/A _09889_/B _09943_/Y vssd1 vssd1 vccd1 vccd1 _09944_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09875_ _13293_/Q vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__inv_2
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08826_ _13653_/Q _08818_/X _08825_/X _08820_/X _08823_/X vssd1 vssd1 vccd1 vccd1
+ _13653_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08757_ _08800_/A vssd1 vssd1 vccd1 vccd1 _08792_/A sky130_fd_sc_hd__buf_4
XPHY_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _07708_/A vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__buf_4
XPHY_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08688_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__buf_2
XPHY_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07639_ _14245_/Q _07634_/X _07313_/X _07636_/X _07624_/X vssd1 vssd1 vccd1 vccd1
+ _14245_/D sky130_fd_sc_hd__o221a_1
XPHY_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _10645_/Y _10425_/X _10646_/Y _10428_/X _10649_/X vssd1 vssd1 vccd1 vccd1
+ _10685_/A sky130_fd_sc_hd__o221a_2
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09309_ _13402_/Q _09302_/X _08146_/A _09303_/X _09306_/X vssd1 vssd1 vccd1 vccd1
+ _13402_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10581_ _10571_/Y _10445_/X _10574_/X _10577_/X _10580_/X vssd1 vssd1 vccd1 vccd1
+ _10603_/C sky130_fd_sc_hd__o2111a_4
XFILLER_126_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12320_ _10340_/Y _14523_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__mux2_4
XFILLER_103_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12251_ _12032_/Y _13352_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11202_ _14619_/Q vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12182_ vssd1 vssd1 vccd1 vccd1 _12182_/HI _12182_/LO sky130_fd_sc_hd__conb_1
XFILLER_135_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11133_ _11131_/Y _10947_/X _11132_/Y _10949_/X vssd1 vssd1 vccd1 vccd1 _11133_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11064_ _14304_/Q vssd1 vssd1 vccd1 vccd1 _11064_/Y sky130_fd_sc_hd__inv_2
XPHY_7030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _13377_/Q _10014_/B _10016_/A vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11966_ _11964_/Y _10195_/A _11965_/Y _10198_/A vssd1 vssd1 vccd1 vccd1 _11966_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ _14183_/CLK _13705_/D vssd1 vssd1 vccd1 vccd1 _13705_/Q sky130_fd_sc_hd__dfxtp_1
X_10917_ _14457_/Q vssd1 vssd1 vccd1 vccd1 _10917_/Y sky130_fd_sc_hd__inv_2
XPHY_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11897_ _14283_/Q vssd1 vssd1 vccd1 vccd1 _11897_/Y sky130_fd_sc_hd__inv_2
XPHY_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ _14146_/CLK _13636_/D vssd1 vssd1 vccd1 vccd1 _13636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10848_ _13949_/Q vssd1 vssd1 vccd1 vccd1 _10848_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ _14120_/CLK _13567_/D vssd1 vssd1 vccd1 vccd1 _13567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10779_ _14337_/Q vssd1 vssd1 vccd1 vccd1 _10779_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12518_ _13366_/Q _10045_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ _14173_/CLK _13498_/D vssd1 vssd1 vccd1 vccd1 _13498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12449_ _12509_/X _06920_/Y _12449_/S vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput505 _12136_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__clkbuf_2
Xoutput516 _12146_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__clkbuf_2
Xoutput527 _12156_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput538 _12166_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput549 _12176_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14119_ _14119_/CLK _14119_/D vssd1 vssd1 vccd1 vccd1 _14119_/Q sky130_fd_sc_hd__dfxtp_1
X_07990_ _14072_/Q _07982_/X _07755_/X _07983_/X _07987_/X vssd1 vssd1 vccd1 vccd1
+ _14072_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06941_ _06954_/A _06941_/B vssd1 vssd1 vccd1 vccd1 _14578_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09660_ _09654_/X _09659_/X _09654_/X _09659_/X vssd1 vssd1 vccd1 vccd1 _09660_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_41_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06872_ _14595_/Q vssd1 vssd1 vccd1 vccd1 _06872_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08611_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08611_/X sky130_fd_sc_hd__buf_1
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09591_ _09597_/A _12337_/X vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__and2_1
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _08554_/A vssd1 vssd1 vccd1 vccd1 _08542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ _08645_/A vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__buf_4
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07424_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07424_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07355_ _14386_/Q _07348_/X _07354_/X _07350_/X _07346_/X vssd1 vssd1 vccd1 vccd1
+ _14386_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ _14415_/Q _07282_/X _06814_/X _07283_/X _07279_/X vssd1 vssd1 vccd1 vccd1
+ _14415_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ _13561_/Q _09022_/X _08933_/X _09023_/X _09019_/X vssd1 vssd1 vccd1 vccd1
+ _13561_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09927_ _09927_/A vssd1 vssd1 vccd1 vccd1 _09927_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09858_ _13310_/Q vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__inv_2
XFILLER_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08809_ _13659_/Q _08748_/A _08577_/X _08750_/A _08808_/X vssd1 vssd1 vccd1 vccd1
+ _13659_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__or2_1
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ _11818_/Y _11693_/X _11819_/Y _11695_/X vssd1 vssd1 vccd1 vccd1 _11820_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_114 _11459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_125 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_158 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _13773_/Q vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__inv_2
XPHY_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_169 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _11412_/A vssd1 vssd1 vccd1 vccd1 _10702_/X sky130_fd_sc_hd__buf_2
XFILLER_202_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14470_ _14470_/CLK _14470_/D vssd1 vssd1 vccd1 vccd1 _14470_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11682_ _14200_/Q vssd1 vssd1 vccd1 vccd1 _11682_/Y sky130_fd_sc_hd__inv_2
XPHY_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13421_ _14173_/CLK _13421_/D vssd1 vssd1 vccd1 vccd1 _13421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10633_ _14178_/Q vssd1 vssd1 vccd1 vccd1 _10633_/Y sky130_fd_sc_hd__inv_2
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13352_ _13352_/CLK _13352_/D vssd1 vssd1 vccd1 vccd1 _13352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10564_ _13663_/Q vssd1 vssd1 vccd1 vccd1 _10564_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _11159_/Y _14540_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13283_ _14538_/CLK _13283_/D vssd1 vssd1 vccd1 vccd1 _13283_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10495_ _11447_/A vssd1 vssd1 vccd1 vccd1 _10495_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12234_/A vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12165_ vssd1 vssd1 vccd1 vccd1 _12165_/HI _12165_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11116_ _11111_/Y _10983_/X _11112_/Y _10985_/X _11115_/X vssd1 vssd1 vccd1 vccd1
+ _11117_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12096_ vssd1 vssd1 vccd1 vccd1 _12096_/HI _12096_/LO sky130_fd_sc_hd__conb_1
XFILLER_42_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11047_ _13875_/Q vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_133_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _12997_/X _12578_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__mux2_1
XPHY_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11949_ _14090_/Q vssd1 vssd1 vccd1 vccd1 _11949_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13619_ _14047_/CLK _13619_/D vssd1 vssd1 vccd1 vccd1 _13619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14599_ _14637_/CLK _14599_/D vssd1 vssd1 vccd1 vccd1 _14599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07140_ _14494_/Q _07136_/X _06810_/X _07137_/X _07139_/X vssd1 vssd1 vccd1 vccd1
+ _14494_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07071_ _07071_/A vssd1 vssd1 vccd1 vccd1 _07071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput368 _12196_/X vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput379 _12197_/X vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07973_ _14082_/Q _07965_/X _07728_/X _07967_/X _07970_/X vssd1 vssd1 vccd1 vccd1
+ _14082_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09712_ _09705_/X _09711_/X _09705_/X _09711_/X vssd1 vssd1 vccd1 vccd1 _10089_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06924_ _14582_/Q vssd1 vssd1 vccd1 vccd1 _06924_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09643_ _14584_/Q _14576_/Q _06915_/Y _06946_/Y vssd1 vssd1 vccd1 vccd1 _09643_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06855_ _09732_/A vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09574_ _09570_/X _09573_/X _13265_/Q _09571_/X vssd1 vssd1 vccd1 vccd1 _13233_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06786_ _14618_/Q _06769_/X _06784_/X _06772_/X _06785_/X vssd1 vssd1 vccd1 vccd1
+ _14618_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08525_ _13804_/Q _08513_/X _08523_/X _08515_/X _08524_/X vssd1 vssd1 vccd1 vccd1
+ _13804_/D sky130_fd_sc_hd__o221a_1
XFILLER_93_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _13835_/Q _08452_/X _08155_/X _08453_/X _08449_/X vssd1 vssd1 vccd1 vccd1
+ _13835_/D sky130_fd_sc_hd__o221a_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07407_ _07484_/A _08340_/B _08584_/C _07630_/D vssd1 vssd1 vccd1 vccd1 _11671_/A
+ sky130_fd_sc_hd__or4_4
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _13872_/Q _08379_/X _08158_/X _08380_/X _08384_/X vssd1 vssd1 vccd1 vccd1
+ _13872_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07338_ _14393_/Q _07335_/X _07336_/X _07337_/X _07333_/X vssd1 vssd1 vccd1 vccd1
+ _14393_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07269_ _14425_/Q _07265_/X _06778_/X _07266_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _14425_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09008_ _13571_/Q _09004_/X _08837_/X _09006_/X _09000_/X vssd1 vssd1 vccd1 vccd1
+ _13571_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10280_ _14327_/Q vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13970_ _14095_/CLK _13970_/D vssd1 vssd1 vccd1 vccd1 _13970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12921_ _12541_/X _12920_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12921_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12524_/X input361/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ _13728_/Q _11642_/X _14047_/Q _11663_/X _11802_/X vssd1 vssd1 vccd1 vccd1
+ _11803_/X sky130_fd_sc_hd__a221o_4
XPHY_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12783_ _09526_/X _12782_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13218_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14637_/CLK _14522_/D vssd1 vssd1 vccd1 vccd1 _14522_/Q sky130_fd_sc_hd__dfxtp_1
X_11734_ _14162_/Q vssd1 vssd1 vccd1 vccd1 _11734_/Y sky130_fd_sc_hd__inv_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11665_ _11665_/A vssd1 vssd1 vccd1 vccd1 _11665_/X sky130_fd_sc_hd__clkbuf_2
X_14453_ _14470_/CLK _14453_/D vssd1 vssd1 vccd1 vccd1 _14453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ _13827_/Q vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13404_ _14188_/CLK _13404_/D vssd1 vssd1 vccd1 vccd1 _13404_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _14627_/CLK _14384_/D vssd1 vssd1 vccd1 vccd1 _14384_/Q sky130_fd_sc_hd__dfxtp_1
X_11596_ _11591_/Y _11397_/X _11592_/Y _11399_/X _11595_/X vssd1 vssd1 vccd1 vccd1
+ _11631_/A sky130_fd_sc_hd__o221a_2
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13352_/CLK _13335_/D vssd1 vssd1 vccd1 vccd1 _13335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10547_ _10542_/Y _10478_/X _10543_/Y _10481_/X _10546_/X vssd1 vssd1 vccd1 vccd1
+ _10560_/B sky130_fd_sc_hd__o221a_4
XFILLER_182_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13266_ _14639_/CLK _13266_/D vssd1 vssd1 vccd1 vccd1 _13266_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10478_ _11435_/A vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12217_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ _14071_/CLK _13197_/D vssd1 vssd1 vccd1 vccd1 _13197_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ vssd1 vssd1 vccd1 vccd1 _12148_/HI _12148_/LO sky130_fd_sc_hd__conb_1
XFILLER_155_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ vssd1 vssd1 vccd1 vccd1 _12079_/HI _12079_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06640_ _08930_/A _06603_/A _06639_/Y _06603_/Y vssd1 vssd1 vccd1 vccd1 _06640_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ _06568_/X _06570_/X _06568_/X _06570_/X vssd1 vssd1 vccd1 vccd1 _06571_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08310_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08310_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09290_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ _13953_/Q _08237_/X _08153_/X _08238_/X _08239_/X vssd1 vssd1 vccd1 vccd1
+ _13953_/D sky130_fd_sc_hd__o221a_1
XANTENNA_14 _11549_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_25 _08217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_36 _08181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _07576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ _08184_/A vssd1 vssd1 vccd1 vccd1 _08172_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_69 _08146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07123_ _14504_/Q _07119_/X _06775_/X _07120_/X _07122_/X vssd1 vssd1 vccd1 vccd1
+ _14504_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07054_ _07071_/A vssd1 vssd1 vccd1 vccd1 _07054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07956_ _08008_/A vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__clkbuf_2
XPHY_6928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06907_ _06901_/X _12295_/X _06906_/Y _06903_/X vssd1 vssd1 vccd1 vccd1 _06908_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07887_ _14129_/Q _07882_/X _07708_/X _07884_/X _07886_/X vssd1 vssd1 vccd1 vccd1
+ _14129_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06838_ _07028_/A vssd1 vssd1 vccd1 vccd1 _06838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ _14567_/Q _09625_/X _14567_/Q _09625_/X vssd1 vssd1 vccd1 vccd1 _09626_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09557_ _09557_/A vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_203_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06769_ _06805_/A vssd1 vssd1 vccd1 vccd1 _06769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08508_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08508_/X sky130_fd_sc_hd__clkbuf_4
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09488_ _13271_/Q _09486_/X _12266_/X _09487_/X vssd1 vssd1 vccd1 vccd1 _13271_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08439_ _13846_/Q _08436_/X _08126_/X _08437_/X _08433_/X vssd1 vssd1 vccd1 vccd1
+ _13846_/D sky130_fd_sc_hd__o221a_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11450_ _14273_/Q vssd1 vssd1 vccd1 vccd1 _11450_/Y sky130_fd_sc_hd__inv_2
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10401_ _13543_/Q _10206_/X _13784_/Q _10209_/X vssd1 vssd1 vccd1 vccd1 _10401_/X
+ sky130_fd_sc_hd__a22o_1
X_11381_ _11376_/Y _11199_/X _11377_/Y _11201_/X _11380_/X vssd1 vssd1 vccd1 vccd1
+ _11394_/B sky130_fd_sc_hd__o221a_1
XFILLER_197_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13120_ _12639_/X input344/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__mux2_1
X_10332_ _10327_/Y _10228_/X _10328_/Y _10231_/X _10331_/X vssd1 vssd1 vccd1 vccd1
+ _10339_/C sky130_fd_sc_hd__o221a_1
XFILLER_137_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13051_ _12604_/X _13050_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10263_ _14210_/Q _10164_/X _14405_/Q _10167_/X _10262_/X vssd1 vssd1 vccd1 vccd1
+ _10298_/B sky130_fd_sc_hd__a221oi_2
XFILLER_69_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12002_ _13857_/Q vssd1 vssd1 vccd1 vccd1 _12002_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10194_ _11658_/A vssd1 vssd1 vccd1 vccd1 _10195_/A sky130_fd_sc_hd__buf_2
XFILLER_94_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13953_ _14107_/CLK _13953_/D vssd1 vssd1 vccd1 vccd1 _13953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _12537_/X input350/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13884_ _14110_/CLK _13884_/D vssd1 vssd1 vccd1 vccd1 _13884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12835_ _12519_/X _12834_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12766_ _09509_/X _12765_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__mux2_1
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14505_ _14621_/CLK _14505_/D vssd1 vssd1 vccd1 vccd1 _14505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11717_ _11715_/Y _11658_/X _11716_/Y _11660_/X vssd1 vssd1 vccd1 vccd1 _11717_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _09597_/X _12696_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _11648_/A vssd1 vssd1 vccd1 vccd1 _11648_/X sky130_fd_sc_hd__clkbuf_2
X_14436_ _14637_/CLK _14436_/D vssd1 vssd1 vccd1 vccd1 _14436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 io_in[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
Xinput23 io_in[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput34 io_in[5] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput45 la_data_in[105] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
XFILLER_50_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14367_ _14633_/CLK _14367_/D vssd1 vssd1 vccd1 vccd1 _14367_/Q sky130_fd_sc_hd__dfxtp_1
X_11579_ _14198_/Q vssd1 vssd1 vccd1 vccd1 _11579_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput56 la_data_in[115] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
XFILLER_171_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput67 la_data_in[125] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_1
Xinput78 la_data_in[1] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_4
XFILLER_116_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput89 la_data_in[2] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__buf_4
X_13318_ _13350_/CLK _13318_/D vssd1 vssd1 vccd1 vccd1 _13318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14298_ _14305_/CLK _14298_/D vssd1 vssd1 vccd1 vccd1 _14298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13249_ _14538_/CLK _13249_/D vssd1 vssd1 vccd1 vccd1 _13281_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08790_ _13671_/Q _08783_/X _08632_/X _08784_/X _08786_/X vssd1 vssd1 vccd1 vccd1
+ _13671_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater613 _12486_/S vssd1 vssd1 vccd1 vccd1 _12603_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater624 _12267_/S vssd1 vssd1 vccd1 vccd1 _12281_/S sky130_fd_sc_hd__buf_8
XFILLER_22_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater635 _13155_/S vssd1 vssd1 vccd1 vccd1 _13179_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07741_ _14195_/Q _07732_/X _07740_/X _07734_/X _07730_/X vssd1 vssd1 vccd1 vccd1
+ _14195_/D sky130_fd_sc_hd__o221a_1
Xrepeater646 _14527_/CLK vssd1 vssd1 vccd1 vccd1 _14611_/CLK sky130_fd_sc_hd__buf_12
Xrepeater657 _14169_/CLK vssd1 vssd1 vccd1 vccd1 _14139_/CLK sky130_fd_sc_hd__buf_12
XFILLER_22_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater668 _14119_/CLK vssd1 vssd1 vccd1 vccd1 _14120_/CLK sky130_fd_sc_hd__buf_12
Xrepeater679 _14071_/CLK vssd1 vssd1 vccd1 vccd1 _14114_/CLK sky130_fd_sc_hd__buf_12
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ _14226_/Q _07669_/X _07365_/X _07670_/X _07666_/X vssd1 vssd1 vccd1 vccd1
+ _14226_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _09413_/A _13059_/X vssd1 vssd1 vccd1 vccd1 _13325_/D sky130_fd_sc_hd__and2_1
X_06623_ _06612_/X _06622_/X _06612_/X _06622_/X vssd1 vssd1 vccd1 vccd1 _06623_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09342_ _09345_/A _12899_/X vssd1 vssd1 vccd1 vccd1 _13381_/D sky130_fd_sc_hd__and2_1
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06554_ _06554_/A vssd1 vssd1 vccd1 vccd1 _06554_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _09327_/A vssd1 vssd1 vccd1 vccd1 _09326_/A sky130_fd_sc_hd__inv_2
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08224_ _13964_/Q _08221_/X _08123_/X _08222_/X _08223_/X vssd1 vssd1 vccd1 vccd1
+ _13964_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08155_ _08155_/A vssd1 vssd1 vccd1 vccd1 _08155_/X sky130_fd_sc_hd__buf_4
XFILLER_181_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07106_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__buf_2
XFILLER_68_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08086_ _14017_/Q _08025_/A _07796_/X _08027_/A _08083_/X vssd1 vssd1 vccd1 vccd1
+ _14017_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ _07130_/A vssd1 vssd1 vccd1 vccd1 _07071_/A sky130_fd_sc_hd__buf_4
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08988_ _13578_/Q _08894_/A _08657_/X _08897_/A _08986_/X vssd1 vssd1 vccd1 vccd1
+ _13578_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07939_ _08133_/A vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__buf_6
XPHY_6758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10950_ _10946_/Y _10947_/X _10948_/Y _10949_/X vssd1 vssd1 vccd1 vccd1 _10950_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09609_ _14587_/Q _14579_/Q _06906_/Y _06933_/Y vssd1 vssd1 vccd1 vccd1 _09610_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_43_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881_ _14067_/Q vssd1 vssd1 vccd1 vccd1 _10881_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _09845_/X _13334_/Q _12650_/S vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ _13290_/Q _12550_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _13487_/Q vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12509_/X _06964_/Y _12482_/S vssd1 vssd1 vccd1 vccd1 _12482_/X sky130_fd_sc_hd__mux2_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11433_ _13216_/Q _11249_/X _14039_/Q _11429_/X _11432_/X vssd1 vssd1 vccd1 vccd1
+ _11433_/X sky130_fd_sc_hd__a221o_4
X_14221_ _14470_/CLK _14221_/D vssd1 vssd1 vccd1 vccd1 _14221_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14152_ _14595_/CLK _14152_/D vssd1 vssd1 vccd1 vccd1 _14152_/Q sky130_fd_sc_hd__dfxtp_1
X_11364_ _13765_/Q vssd1 vssd1 vccd1 vccd1 _11364_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10315_ _13977_/Q vssd1 vssd1 vccd1 vccd1 _10315_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _12629_/X _13102_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14083_ _14291_/CLK _14083_/D vssd1 vssd1 vccd1 vccd1 _14083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11295_ _14348_/Q vssd1 vssd1 vccd1 vccd1 _11295_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13034_ _13033_/X _12596_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13034_/X sky130_fd_sc_hd__mux2_1
X_10246_ _13461_/Q vssd1 vssd1 vccd1 vccd1 _10246_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10177_ _11646_/A vssd1 vssd1 vccd1 vccd1 _10178_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13936_ _14095_/CLK _13936_/D vssd1 vssd1 vccd1 vccd1 _13936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13867_ _14107_/CLK _13867_/D vssd1 vssd1 vccd1 vccd1 _13867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ _12516_/X _12817_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12818_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13798_ _14114_/CLK _13798_/D vssd1 vssd1 vccd1 vccd1 _13798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _09550_/X _12748_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14419_ _14538_/CLK _14419_/D vssd1 vssd1 vccd1 vccd1 _14419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09960_ _13291_/Q _09958_/Y _09886_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08911_ _13609_/Q _08905_/X _08606_/X _08907_/X _08910_/X vssd1 vssd1 vccd1 vccd1
+ _13609_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__or2_1
XFILLER_174_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08842_ _13647_/Q _08832_/X _08508_/X _08835_/X _08839_/X vssd1 vssd1 vccd1 vccd1
+ _13647_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08773_ _13681_/Q _08767_/X _08521_/X _08768_/X _08769_/X vssd1 vssd1 vccd1 vccd1
+ _13681_/D sky130_fd_sc_hd__o221a_1
XPHY_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07724_ _14202_/Q _07718_/X _07723_/X _07721_/X _07715_/X vssd1 vssd1 vccd1 vccd1
+ _14202_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07655_ _14237_/Q _07653_/X _07336_/X _07654_/X _07650_/X vssd1 vssd1 vccd1 vccd1
+ _14237_/D sky130_fd_sc_hd__o221a_1
XPHY_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06606_ _06592_/X _06605_/X _06592_/X _06605_/X vssd1 vssd1 vccd1 vccd1 _06606_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07586_ _14274_/Q _07580_/X _07341_/X _07581_/X _07585_/X vssd1 vssd1 vccd1 vccd1
+ _14274_/D sky130_fd_sc_hd__o221a_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09325_ _13392_/Q _09318_/X _08171_/A _09319_/X _09322_/X vssd1 vssd1 vccd1 vccd1
+ _13392_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06537_ _08833_/A _08837_/A _06535_/Y _06536_/Y vssd1 vssd1 vccd1 vccd1 _06537_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _13431_/Q _09249_/X _08967_/X _09250_/X _09252_/X vssd1 vssd1 vccd1 vccd1
+ _13431_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ _13972_/Q _08198_/X _08101_/X _08201_/X _08204_/X vssd1 vssd1 vccd1 vccd1
+ _13972_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09187_ _13470_/Q _09179_/X _08967_/X _09180_/X _09182_/X vssd1 vssd1 vccd1 vccd1
+ _13470_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08138_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08069_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10100_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__buf_2
XFILLER_1_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11080_ _13674_/Q vssd1 vssd1 vccd1 vccd1 _11080_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _13368_/Q _09994_/B _09995_/A vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__o21a_1
Xinput202 la_oenb[16] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_1
XFILLER_66_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput213 la_oenb[26] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_1
XFILLER_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput224 la_oenb[36] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_1
XPHY_7245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 la_oenb[46] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_1
XPHY_7256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput246 la_oenb[56] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_1
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput257 la_oenb[66] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__buf_1
XFILLER_44_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput268 la_oenb[76] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__buf_1
XPHY_7289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput279 la_oenb[86] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_hd__buf_1
XFILLER_40_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _13934_/Q vssd1 vssd1 vccd1 vccd1 _11982_/Y sky130_fd_sc_hd__inv_2
XPHY_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13721_ _14143_/CLK _13721_/D vssd1 vssd1 vccd1 vccd1 _13721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10933_ _11406_/A vssd1 vssd1 vccd1 vccd1 _10933_/X sky130_fd_sc_hd__clkbuf_4
XPHY_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13652_ _14056_/CLK _13652_/D vssd1 vssd1 vccd1 vccd1 _13652_/Q sky130_fd_sc_hd__dfxtp_1
X_10864_ _14378_/Q vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _09907_/Y _13311_/Q _12603_/S vssd1 vssd1 vccd1 vccd1 _12603_/X sky130_fd_sc_hd__mux2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _14178_/CLK _13583_/D vssd1 vssd1 vccd1 vccd1 _13583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10790_/Y _10745_/X _10791_/Y _10747_/X _10794_/X vssd1 vssd1 vccd1 vccd1
+ _10796_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12534_ _13382_/Q _10029_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12534_/X sky130_fd_sc_hd__mux2_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12465_ _12464_/X _06938_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12465_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204_ _14325_/CLK _14204_/D vssd1 vssd1 vccd1 vccd1 _14204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11416_ _11416_/A vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12396_ _13222_/Q _12395_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _14139_/CLK _14135_/D vssd1 vssd1 vccd1 vccd1 _14135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11347_ _13920_/Q vssd1 vssd1 vccd1 vccd1 _11347_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ _11514_/A vssd1 vssd1 vccd1 vccd1 _11278_/X sky130_fd_sc_hd__buf_2
XFILLER_106_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14066_ _14143_/CLK _14066_/D vssd1 vssd1 vccd1 vccd1 _14066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10229_ _13578_/Q vssd1 vssd1 vccd1 vccd1 _10229_/Y sky130_fd_sc_hd__inv_2
X_13017_ _12588_/X _13016_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13919_ _14146_/CLK _13919_/D vssd1 vssd1 vccd1 vccd1 _13919_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07440_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07440_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07371_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07371_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _13514_/Q _09103_/X _08954_/X _09104_/X _09109_/X vssd1 vssd1 vccd1 vccd1
+ _13514_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09041_ _13552_/Q _09039_/X _08957_/X _09040_/X _09036_/X vssd1 vssd1 vccd1 vccd1
+ _13552_/D sky130_fd_sc_hd__o221a_1
Xclkbuf_2_3_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _13350_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_148_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09943_ _09943_/A vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09874_ _13294_/Q vssd1 vssd1 vccd1 vccd1 _09888_/A sky130_fd_sc_hd__inv_2
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08825_ _08825_/A vssd1 vssd1 vccd1 vccd1 _08825_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _13690_/Q _08748_/X _08496_/X _08750_/X _08751_/X vssd1 vssd1 vccd1 vccd1
+ _13690_/D sky130_fd_sc_hd__o221a_1
XPHY_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07707_ _14208_/Q _07704_/X _07412_/X _07706_/X _07698_/X vssd1 vssd1 vccd1 vccd1
+ _14208_/D sky130_fd_sc_hd__o221a_1
XPHY_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08687_/X sky130_fd_sc_hd__buf_2
XPHY_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07638_ _14246_/Q _07634_/X _07311_/X _07636_/X _07624_/X vssd1 vssd1 vccd1 vccd1
+ _14246_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07569_ _14282_/Q _07561_/X _07317_/X _07563_/X _07566_/X vssd1 vssd1 vccd1 vccd1
+ _14282_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09308_ _13403_/Q _09302_/X _08144_/A _09303_/X _09306_/X vssd1 vssd1 vccd1 vccd1
+ _13403_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10580_ _10578_/Y _10462_/X _10579_/Y _10465_/X vssd1 vssd1 vccd1 vccd1 _10580_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ _13442_/Q _09233_/X _08940_/X _09234_/X _09236_/X vssd1 vssd1 vccd1 vccd1
+ _13442_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _12031_/Y _13351_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12250_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11201_ _11437_/A vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12181_ vssd1 vssd1 vccd1 vccd1 _12181_/HI _12181_/LO sky130_fd_sc_hd__conb_1
XFILLER_162_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11132_ _14111_/Q vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11063_ _11058_/Y _10963_/X _11059_/Y _10965_/X _11062_/X vssd1 vssd1 vccd1 vccd1
+ _11076_/B sky130_fd_sc_hd__o221a_4
XPHY_7020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _13377_/Q _10014_/B vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11965_ _13537_/Q vssd1 vssd1 vccd1 vccd1 _11965_/Y sky130_fd_sc_hd__inv_2
XPHY_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _14183_/CLK _13704_/D vssd1 vssd1 vccd1 vccd1 _13704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10916_ _13475_/Q vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11896_ _14205_/Q vssd1 vssd1 vccd1 vccd1 _11896_/Y sky130_fd_sc_hd__inv_2
XPHY_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13635_ _14071_/CLK _13635_/D vssd1 vssd1 vccd1 vccd1 _13635_/Q sky130_fd_sc_hd__dfxtp_1
X_10847_ _14222_/Q _10696_/X _14417_/Q _10697_/X _10846_/X vssd1 vssd1 vccd1 vccd1
+ _10880_/B sky130_fd_sc_hd__a221oi_2
XFILLER_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13566_ _14120_/CLK _13566_/D vssd1 vssd1 vccd1 vccd1 _13566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10778_ _14493_/Q vssd1 vssd1 vccd1 vccd1 _10778_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _13352_/Q _10049_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12517_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13497_ _14173_/CLK _13497_/D vssd1 vssd1 vccd1 vccd1 _13497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _12447_/X _06915_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput506 _12137_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput517 _12147_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput528 _12157_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput539 _12167_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__clkbuf_2
X_12379_ _12378_/X _13212_/Q _12645_/S vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14118_ _14119_/CLK _14118_/D vssd1 vssd1 vccd1 vccd1 _14118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06940_ _06937_/X _12304_/X _06938_/Y _06939_/X vssd1 vssd1 vccd1 vccd1 _06941_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14049_ _14056_/CLK _14049_/D vssd1 vssd1 vccd1 vccd1 _14049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06871_ _06877_/A _06871_/B vssd1 vssd1 vccd1 vccd1 _14596_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08610_ _08635_/A vssd1 vssd1 vccd1 vccd1 _08610_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09590_ _09583_/X _09589_/X _13259_/Q _09584_/X vssd1 vssd1 vccd1 vccd1 _13227_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08541_ _08945_/A vssd1 vssd1 vccd1 vccd1 _08541_/X sky130_fd_sc_hd__buf_4
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08472_ _13825_/Q _08468_/X _08179_/X _08469_/X _08465_/X vssd1 vssd1 vccd1 vccd1
+ _13825_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07423_ _07468_/A vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _08142_/A vssd1 vssd1 vccd1 vccd1 _07354_/X sky130_fd_sc_hd__buf_2
XFILLER_52_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07285_ _14416_/Q _07282_/X _06810_/X _07283_/X _07279_/X vssd1 vssd1 vccd1 vccd1
+ _14416_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09024_ _13562_/Q _09022_/X _08930_/X _09023_/X _09019_/X vssd1 vssd1 vccd1 vccd1
+ _13562_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09926_ _09926_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__or2_1
XFILLER_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09857_ _13311_/Q vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__inv_2
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08808_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09788_ _09788_/A _09824_/A vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__or2_2
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _13698_/Q _08677_/A _08577_/X _08679_/A _08737_/X vssd1 vssd1 vccd1 vccd1
+ _13698_/D sky130_fd_sc_hd__o221a_1
XPHY_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _09545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_115 _11461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_137 _11359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11750_ _13968_/Q vssd1 vssd1 vccd1 vccd1 _11750_/Y sky130_fd_sc_hd__inv_2
XPHY_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _11947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _13946_/Q vssd1 vssd1 vccd1 vccd1 _10701_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A vssd1 vssd1 vccd1 vccd1 _11681_/X sky130_fd_sc_hd__buf_2
XPHY_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _14173_/CLK _13420_/D vssd1 vssd1 vccd1 vccd1 _13420_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _13586_/Q vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__inv_2
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10563_ _13429_/Q vssd1 vssd1 vccd1 vccd1 _10563_/Y sky130_fd_sc_hd__inv_2
X_13351_ _13370_/CLK _13351_/D vssd1 vssd1 vccd1 vccd1 _13351_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _11229_/Y _14541_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__mux2_1
X_10494_ _11681_/A vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__buf_4
X_13282_ _14538_/CLK _13282_/D vssd1 vssd1 vccd1 vccd1 _13282_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12233_ _12233_/A vssd1 vssd1 vccd1 vccd1 _12233_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12164_ vssd1 vssd1 vccd1 vccd1 _12164_/HI _12164_/LO sky130_fd_sc_hd__conb_1
XFILLER_194_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11115_ _11113_/Y _10987_/X _11114_/Y _10989_/X vssd1 vssd1 vccd1 vccd1 _11115_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ vssd1 vssd1 vccd1 vccd1 _12095_/HI _12095_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11046_ _13758_/Q vssd1 vssd1 vccd1 vccd1 _11046_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _12578_/X _12996_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ _11948_/A _11948_/B _11948_/C _11948_/D vssd1 vssd1 vccd1 vccd1 _11948_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_166_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ _13854_/Q vssd1 vssd1 vccd1 vccd1 _11879_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13618_ _14047_/CLK _13618_/D vssd1 vssd1 vccd1 vccd1 _13618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14598_ _14621_/CLK _14598_/D vssd1 vssd1 vccd1 vccd1 _14598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13549_ _14120_/CLK _13549_/D vssd1 vssd1 vccd1 vccd1 _13549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07070_ _07070_/A vssd1 vssd1 vccd1 vccd1 _07070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput369 _12206_/X vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07972_ _14083_/Q _07965_/X _07726_/X _07967_/X _07970_/X vssd1 vssd1 vccd1 vccd1
+ _14083_/D sky130_fd_sc_hd__o221a_1
XFILLER_155_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09711_ _09706_/X _09710_/X _09706_/X _09710_/X vssd1 vssd1 vccd1 vccd1 _09711_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06923_ _06935_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _14583_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09642_ _09640_/A _09641_/A _09640_/Y _09641_/Y vssd1 vssd1 vccd1 vccd1 _09642_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06854_ _06918_/A vssd1 vssd1 vccd1 vccd1 _06877_/A sky130_fd_sc_hd__buf_1
XFILLER_186_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09573_/A _12364_/X vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__and2_1
X_06785_ _06785_/A vssd1 vssd1 vccd1 vccd1 _06785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08524_ _08524_/A vssd1 vssd1 vccd1 vccd1 _08524_/X sky130_fd_sc_hd__buf_2
XFILLER_97_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ _13836_/Q _08452_/X _08153_/X _08453_/X _08449_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07406_ _08482_/B vssd1 vssd1 vccd1 vccd1 _08340_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ _13873_/Q _08379_/X _08243_/X _08380_/X _08384_/X vssd1 vssd1 vccd1 vccd1
+ _13873_/D sky130_fd_sc_hd__o221a_1
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07337_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07268_ _14426_/Q _07265_/X _06775_/X _07266_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _14426_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09007_ _13572_/Q _09004_/X _08833_/X _09006_/X _09000_/X vssd1 vssd1 vccd1 vccd1
+ _13572_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07199_ _14463_/Q _07193_/X _06781_/X _07194_/X _07197_/X vssd1 vssd1 vccd1 vccd1
+ _14463_/D sky130_fd_sc_hd__o221a_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09909_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__or2_2
XFILLER_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12920_ _12541_/X input346/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12851_ _12523_/X _12850_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__mux2_1
XPHY_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11802_ _13572_/Q _11664_/X _13813_/Q _11665_/X vssd1 vssd1 vccd1 vccd1 _11802_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _09526_/X _12781_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14521_ _14637_/CLK _14521_/D vssd1 vssd1 vccd1 vccd1 _14521_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _13928_/Q vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__inv_2
XPHY_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14452_ _14470_/CLK _14452_/D vssd1 vssd1 vccd1 vccd1 _14452_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _14188_/CLK _13403_/D vssd1 vssd1 vccd1 vccd1 _13403_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10615_ _10613_/Y _10448_/X _10614_/Y _10451_/X vssd1 vssd1 vccd1 vccd1 _10615_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14383_ _14627_/CLK _14383_/D vssd1 vssd1 vccd1 vccd1 _14383_/Q sky130_fd_sc_hd__dfxtp_1
X_11595_ _11593_/Y _11401_/X _11594_/Y _11403_/X vssd1 vssd1 vccd1 vccd1 _11595_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13334_ _13352_/CLK _13334_/D vssd1 vssd1 vccd1 vccd1 _13334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10546_ _10544_/Y _10484_/X _10545_/Y _10487_/X vssd1 vssd1 vccd1 vccd1 _10546_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _14639_/CLK _13265_/D vssd1 vssd1 vccd1 vccd1 _13265_/Q sky130_fd_sc_hd__dfxtp_2
X_10477_ _11669_/A vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__buf_2
XFILLER_124_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12216_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13196_ _14071_/CLK _13196_/D vssd1 vssd1 vccd1 vccd1 _13196_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12147_ vssd1 vssd1 vccd1 vccd1 _12147_/HI _12147_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12078_ vssd1 vssd1 vccd1 vccd1 _12078_/HI _12078_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11029_ _14147_/Q vssd1 vssd1 vccd1 vccd1 _11029_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _08945_/A _06556_/Y _06569_/Y _08954_/A vssd1 vssd1 vccd1 vccd1 _06570_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08240_ _13954_/Q _08237_/X _08150_/X _08238_/X _08239_/X vssd1 vssd1 vccd1 vccd1
+ _13954_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_15 _11699_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_26 _08217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_37 _06843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08171_ _08171_/A vssd1 vssd1 vccd1 vccd1 _08171_/X sky130_fd_sc_hd__buf_4
XANTENNA_48 _07679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_59 _07788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ _07062_/A vssd1 vssd1 vccd1 vccd1 _07053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ _07955_/A vssd1 vssd1 vccd1 vccd1 _07955_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06906_ _14587_/Q vssd1 vssd1 vccd1 vccd1 _06906_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07886_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__buf_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09625_ _06865_/X _09624_/X _06865_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _09625_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06837_ _08183_/A vssd1 vssd1 vccd1 vccd1 _06837_/X sky130_fd_sc_hd__buf_2
XFILLER_186_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _09560_/A _12394_/X vssd1 vssd1 vccd1 vccd1 _09556_/X sky130_fd_sc_hd__and2_1
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06768_ _14623_/Q _06751_/X _06766_/X _06754_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _14623_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08507_ _13811_/Q _08500_/X _08217_/X _08503_/X _08497_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/D sky130_fd_sc_hd__o221a_1
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09487_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09487_/X sky130_fd_sc_hd__clkbuf_2
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06699_ _06699_/A vssd1 vssd1 vccd1 vccd1 _06699_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08438_ _13847_/Q _08436_/X _08123_/X _08437_/X _08433_/X vssd1 vssd1 vccd1 vccd1
+ _13847_/D sky130_fd_sc_hd__o221a_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08369_ _13883_/Q _08363_/X _08130_/X _08364_/X _08367_/X vssd1 vssd1 vccd1 vccd1
+ _13883_/D sky130_fd_sc_hd__o221a_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10400_ _10390_/Y _10178_/X _10393_/X _10396_/X _10399_/X vssd1 vssd1 vccd1 vccd1
+ _10422_/C sky130_fd_sc_hd__o2111a_4
XFILLER_109_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11380_ _11378_/Y _11203_/X _11379_/Y _11205_/X vssd1 vssd1 vccd1 vccd1 _11380_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _10329_/Y _10234_/X _10330_/Y _10237_/X vssd1 vssd1 vccd1 vccd1 _10331_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10262_ _13384_/Q _11747_/A _13696_/Q _10173_/X vssd1 vssd1 vccd1 vccd1 _10262_/X
+ sky130_fd_sc_hd__a22o_1
X_13050_ _13049_/X _12604_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13050_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12001_ _11999_/Y _10181_/A _12000_/Y _10184_/A vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _13975_/Q vssd1 vssd1 vccd1 vccd1 _10193_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13952_ _14107_/CLK _13952_/D vssd1 vssd1 vccd1 vccd1 _13952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12903_ _12536_/X _12902_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12903_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13883_ _14110_/CLK _13883_/D vssd1 vssd1 vccd1 vccd1 _13883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12834_ _12519_/X _12833_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12834_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12765_ _09509_/X _12764_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14504_ _14621_/CLK _14504_/D vssd1 vssd1 vccd1 vccd1 _14504_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _13531_/Q vssd1 vssd1 vccd1 vccd1 _11716_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12696_ _09597_/X input330/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__mux2_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14435_ _14527_/CLK _14435_/D vssd1 vssd1 vccd1 vccd1 _14435_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _13771_/Q vssd1 vssd1 vccd1 vccd1 _11647_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 io_in[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_141_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput24 io_in[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
Xinput35 io_in[6] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
X_14366_ _14633_/CLK _14366_/D vssd1 vssd1 vccd1 vccd1 _14366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11578_ _13606_/Q vssd1 vssd1 vccd1 vccd1 _11578_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput46 la_data_in[106] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
XFILLER_200_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput57 la_data_in[116] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 la_data_in[126] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_1
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13317_ _14459_/CLK _13317_/D vssd1 vssd1 vccd1 vccd1 _13317_/Q sky130_fd_sc_hd__dfxtp_1
X_10529_ _13747_/Q vssd1 vssd1 vccd1 vccd1 _10529_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput79 la_data_in[20] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_1
X_14297_ _14305_/CLK _14297_/D vssd1 vssd1 vccd1 vccd1 _14297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _13350_/CLK _13248_/D vssd1 vssd1 vccd1 vccd1 _13280_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13179_ _12667_/X _13178_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater614 _13146_/S vssd1 vssd1 vccd1 vccd1 _13178_/S sky130_fd_sc_hd__buf_8
XFILLER_26_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater625 _12262_/S vssd1 vssd1 vccd1 vccd1 _12267_/S sky130_fd_sc_hd__buf_6
XFILLER_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ _08130_/A vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__buf_4
XFILLER_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater636 _13147_/S vssd1 vssd1 vccd1 vccd1 _13155_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_61_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater647 _14633_/CLK vssd1 vssd1 vccd1 vccd1 _14629_/CLK sky130_fd_sc_hd__buf_12
XFILLER_26_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater658 _14169_/CLK vssd1 vssd1 vccd1 vccd1 _14173_/CLK sky130_fd_sc_hd__buf_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater669 _14183_/CLK vssd1 vssd1 vccd1 vccd1 _14188_/CLK sky130_fd_sc_hd__buf_12
XFILLER_93_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _14227_/Q _07669_/X _07362_/X _07670_/X _07666_/X vssd1 vssd1 vccd1 vccd1
+ _14227_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09410_ _09413_/A _13055_/X vssd1 vssd1 vccd1 vccd1 _13326_/D sky130_fd_sc_hd__and2_1
XFILLER_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06622_ _06615_/X _06621_/X _06615_/X _06621_/X vssd1 vssd1 vccd1 vccd1 _06622_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09341_ _09345_/A _12895_/X vssd1 vssd1 vccd1 vccd1 _13382_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06553_ _06553_/A vssd1 vssd1 vccd1 vccd1 _06553_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09272_ _09272_/A _10168_/A vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__or2_2
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08223_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08154_ _13992_/Q _08149_/X _08153_/X _08151_/X _08147_/X vssd1 vssd1 vccd1 vccd1
+ _13992_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07105_ _14515_/Q _07102_/X _06735_/X _07104_/X _07096_/X vssd1 vssd1 vccd1 vccd1
+ _14515_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08085_ _14018_/Q _08078_/X _07792_/X _08079_/X _08083_/X vssd1 vssd1 vccd1 vccd1
+ _14018_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07036_ _07062_/A vssd1 vssd1 vccd1 vccd1 _07036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _13579_/Q _08894_/A _08985_/X _08897_/A _08986_/X vssd1 vssd1 vccd1 vccd1
+ _13579_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__buf_2
XFILLER_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07869_ _14137_/Q _07863_/X _07788_/X _07864_/X _07865_/X vssd1 vssd1 vccd1 vccd1
+ _14137_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _06952_/Y _14570_/Q _14574_/Q _06967_/Y vssd1 vssd1 vccd1 vccd1 _09608_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _10880_/A _10880_/B _10880_/C _10880_/D vssd1 vssd1 vccd1 vccd1 _10880_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_186_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _09547_/A _12373_/X vssd1 vssd1 vccd1 vccd1 _09539_/X sky130_fd_sc_hd__and2_1
XFILLER_38_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ _09959_/Y _13290_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _14157_/Q vssd1 vssd1 vccd1 vccd1 _11501_/Y sky130_fd_sc_hd__inv_2
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12480_/X _06961_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12481_/X sky130_fd_sc_hd__mux2_2
XFILLER_40_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14220_ _14470_/CLK _14220_/D vssd1 vssd1 vccd1 vccd1 _14220_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _13564_/Q _11430_/X _13805_/Q _11431_/X vssd1 vssd1 vccd1 vccd1 _11432_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14305_/CLK _14151_/D vssd1 vssd1 vccd1 vccd1 _14151_/Q sky130_fd_sc_hd__dfxtp_1
X_11363_ _13960_/Q vssd1 vssd1 vccd1 vccd1 _11363_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _13101_/X _12629_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__mux2_1
X_10314_ _10312_/Y _10188_/X _10313_/Y _10191_/X vssd1 vssd1 vccd1 vccd1 _10314_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14082_ _14291_/CLK _14082_/D vssd1 vssd1 vccd1 vccd1 _14082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11294_ _14504_/Q vssd1 vssd1 vccd1 vccd1 _11294_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ _12596_/X _13032_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _13033_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10245_ _10245_/A vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10176_ _13936_/Q vssd1 vssd1 vccd1 vccd1 _10176_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13935_ _14169_/CLK _13935_/D vssd1 vssd1 vccd1 vccd1 _13935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13866_ _14100_/CLK _13866_/D vssd1 vssd1 vccd1 vccd1 _13866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12817_ _12516_/X _12816_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13797_ _14114_/CLK _13797_/D vssd1 vssd1 vccd1 vccd1 _13797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12748_ _09550_/X input340/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12679_ _09586_/X _12678_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13196_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14418_ _14538_/CLK _14418_/D vssd1 vssd1 vccd1 vccd1 _14418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14349_ _14627_/CLK _14349_/D vssd1 vssd1 vccd1 vccd1 _14349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08910_ _08923_/A vssd1 vssd1 vccd1 vccd1 _08910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09890_ _09890_/A _09943_/A vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__or2_1
XFILLER_48_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08841_ _13648_/Q _08832_/X _08606_/X _08835_/X _08839_/X vssd1 vssd1 vccd1 vccd1
+ _13648_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08772_ _13682_/Q _08767_/X _08519_/X _08768_/X _08769_/X vssd1 vssd1 vccd1 vccd1
+ _13682_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07723_ _07723_/A vssd1 vssd1 vccd1 vccd1 _07723_/X sky130_fd_sc_hd__buf_4
XFILLER_187_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07654_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07654_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06605_ _06599_/X _06604_/X _06599_/X _06604_/X vssd1 vssd1 vccd1 vccd1 _06605_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07585_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07585_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _13393_/Q _09318_/X _08169_/A _09319_/X _09322_/X vssd1 vssd1 vccd1 vccd1
+ _13393_/D sky130_fd_sc_hd__o221a_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06536_ _06536_/A vssd1 vssd1 vccd1 vccd1 _06536_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _13432_/Q _09249_/X _08965_/X _09250_/X _09252_/X vssd1 vssd1 vccd1 vccd1
+ _13432_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08206_ _13973_/Q _08198_/X _08099_/X _08201_/X _08204_/X vssd1 vssd1 vccd1 vccd1
+ _13973_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09186_ _13471_/Q _09179_/X _08965_/X _09180_/X _09182_/X vssd1 vssd1 vccd1 vccd1
+ _13471_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08137_ _08137_/A vssd1 vssd1 vccd1 vccd1 _08137_/X sky130_fd_sc_hd__buf_4
XFILLER_134_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ _14028_/Q _08061_/X _07767_/X _08062_/X _08066_/X vssd1 vssd1 vccd1 vccd1
+ _14028_/D sky130_fd_sc_hd__o221a_1
XFILLER_150_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07019_ _14559_/Q _07014_/X _07015_/X _07017_/X _07018_/X vssd1 vssd1 vccd1 vccd1
+ _14559_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10030_ _13367_/Q _09992_/B _09993_/A vssd1 vssd1 vccd1 vccd1 _10030_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput203 la_oenb[17] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__buf_1
XPHY_7224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 la_oenb[27] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__buf_1
XPHY_7235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput225 la_oenb[37] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_1
XFILLER_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput236 la_oenb[47] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_1
XPHY_7257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput247 la_oenb[57] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__buf_1
XPHY_7268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 la_oenb[67] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__buf_1
XFILLER_44_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput269 la_oenb[77] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__buf_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _11976_/Y _10228_/A _11977_/Y _10231_/A _11980_/X vssd1 vssd1 vccd1 vccd1
+ _11988_/C sky130_fd_sc_hd__o221a_1
XPHY_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13720_ _14183_/CLK _13720_/D vssd1 vssd1 vccd1 vccd1 _13720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10932_ _11830_/A vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__buf_4
XFILLER_79_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _14056_/CLK _13651_/D vssd1 vssd1 vccd1 vccd1 _13651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10863_ _14612_/Q vssd1 vssd1 vccd1 vccd1 _10863_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _13312_/Q _12601_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13582_ _14178_/CLK _13582_/D vssd1 vssd1 vccd1 vccd1 _13582_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _10792_/Y _10749_/X _10793_/Y _10751_/X vssd1 vssd1 vccd1 vccd1 _10794_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ _13367_/Q _10030_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12464_ _12509_/X _06938_/Y _12464_/S vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14203_ _14481_/CLK _14203_/D vssd1 vssd1 vccd1 vccd1 _14203_/Q sky130_fd_sc_hd__dfxtp_1
X_11415_ _13883_/Q vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ _13222_/Q _06743_/Y _12407_/S vssd1 vssd1 vccd1 vccd1 _12395_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _14173_/CLK _14134_/D vssd1 vssd1 vccd1 vccd1 _14134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _11341_/Y _11209_/X _11342_/Y _11211_/X _11345_/X vssd1 vssd1 vccd1 vccd1
+ _11353_/C sky130_fd_sc_hd__o221a_1
XFILLER_173_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14065_ _14143_/CLK _14065_/D vssd1 vssd1 vccd1 vccd1 _14065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11277_ _11272_/Y _11161_/X _11273_/Y _11163_/X _11276_/X vssd1 vssd1 vccd1 vccd1
+ _11313_/A sky130_fd_sc_hd__o221a_2
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ _12588_/X input337/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10228_ _10228_/A vssd1 vssd1 vccd1 vccd1 _10228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10159_ _10159_/A vssd1 vssd1 vccd1 vccd1 _10159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918_ _14146_/CLK _13918_/D vssd1 vssd1 vccd1 vccd1 _13918_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13849_ _14094_/CLK _13849_/D vssd1 vssd1 vccd1 vccd1 _13849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ _08158_/A vssd1 vssd1 vccd1 vccd1 _07370_/X sky130_fd_sc_hd__buf_4
XFILLER_17_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09040_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09942_ _13310_/Q _09940_/Y _09905_/B vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09873_ _13295_/Q vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__inv_2
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08824_ _13654_/Q _08818_/X _08822_/X _08820_/X _08823_/X vssd1 vssd1 vccd1 vccd1
+ _13654_/D sky130_fd_sc_hd__o221a_1
XFILLER_86_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _13691_/Q _08748_/X _08494_/X _08750_/X _08751_/X vssd1 vssd1 vccd1 vccd1
+ _13691_/D sky130_fd_sc_hd__o221a_1
XPHY_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07706_ _07706_/A vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08686_ _08730_/A vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__buf_2
XPHY_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07637_ _14247_/Q _07634_/X _07412_/X _07636_/X _07624_/X vssd1 vssd1 vccd1 vccd1
+ _14247_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07568_ _14283_/Q _07561_/X _07315_/X _07563_/X _07566_/X vssd1 vssd1 vccd1 vccd1
+ _14283_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09307_ _13404_/Q _09302_/X _08142_/A _09303_/X _09306_/X vssd1 vssd1 vccd1 vccd1
+ _13404_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06519_ _08813_/A vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__buf_2
XFILLER_167_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07499_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _13443_/Q _09233_/X _08935_/X _09234_/X _09236_/X vssd1 vssd1 vccd1 vccd1
+ _13443_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09169_ _13481_/Q _09163_/X _08940_/X _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1
+ _13481_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11200_ _14346_/Q vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12180_ vssd1 vssd1 vccd1 vccd1 _12180_/HI _12180_/LO sky130_fd_sc_hd__conb_1
XFILLER_194_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _13838_/Q vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11062_ _11060_/Y _10967_/X _11061_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _11062_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10013_ _10013_/A vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__inv_2
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _14012_/Q vssd1 vssd1 vccd1 vccd1 _11964_/Y sky130_fd_sc_hd__inv_2
XPHY_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _14178_/CLK _13703_/D vssd1 vssd1 vccd1 vccd1 _13703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10915_ _14145_/Q vssd1 vssd1 vccd1 vccd1 _10915_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11895_ _13613_/Q vssd1 vssd1 vccd1 vccd1 _11895_/Y sky130_fd_sc_hd__inv_2
XPHY_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13634_ _14071_/CLK _13634_/D vssd1 vssd1 vccd1 vccd1 _13634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10846_ _13396_/Q _10804_/X _13708_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _10846_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13565_ _14120_/CLK _13565_/D vssd1 vssd1 vccd1 vccd1 _13565_/Q sky130_fd_sc_hd__dfxtp_1
X_10777_ _13202_/Q _10775_/X _14025_/Q _10719_/X _10776_/X vssd1 vssd1 vccd1 vccd1
+ _10777_/X sky130_fd_sc_hd__a221o_2
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12516_ _13353_/Q _10050_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12516_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13496_ _14173_/CLK _13496_/D vssd1 vssd1 vccd1 vccd1 _13496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12447_ _12446_/X _06915_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12447_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput507 _12138_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput518 _12148_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12378_ _13212_/Q _12377_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput529 _12158_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14117_ _14119_/CLK _14117_/D vssd1 vssd1 vccd1 vccd1 _14117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11329_ _13998_/Q vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14048_ _14056_/CLK _14048_/D vssd1 vssd1 vccd1 vccd1 _14048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06870_ _06857_/X _12286_/X _06869_/X _06861_/X vssd1 vssd1 vccd1 vccd1 _06871_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08540_ _08552_/A vssd1 vssd1 vccd1 vccd1 _08540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08471_ _13826_/Q _08468_/X _08259_/X _08469_/X _08465_/X vssd1 vssd1 vccd1 vccd1
+ _13826_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07422_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07353_ _14387_/Q _07348_/X _07352_/X _07350_/X _07346_/X vssd1 vssd1 vccd1 vccd1
+ _14387_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07284_ _14417_/Q _07282_/X _06807_/X _07283_/X _07279_/X vssd1 vssd1 vccd1 vccd1
+ _14417_/D sky130_fd_sc_hd__o221a_1
XFILLER_176_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09023_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09925_ _13317_/Q vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__inv_2
XFILLER_28_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09856_ _09776_/A _09776_/B _09777_/B vssd1 vssd1 vccd1 vccd1 _09856_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_115_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08807_ _13660_/Q _08800_/X _08574_/X _08801_/X _08802_/X vssd1 vssd1 vccd1 vccd1
+ _13660_/D sky130_fd_sc_hd__o221a_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ _09787_/A _09787_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__or2_2
XFILLER_22_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06999_ _14561_/Q vssd1 vssd1 vccd1 vccd1 _06999_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08738_ _13699_/Q _08730_/X _08574_/X _08731_/X _08737_/X vssd1 vssd1 vccd1 vccd1
+ _13699_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_116 _10541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _11375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08669_ _13736_/Q _08662_/X _08496_/X _08663_/X _08665_/X vssd1 vssd1 vccd1 vccd1
+ _13736_/D sky130_fd_sc_hd__o221a_1
XANTENNA_149 _11500_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10700_ _14219_/Q _10696_/X _14414_/Q _10697_/X _10699_/X vssd1 vssd1 vccd1 vccd1
+ _10755_/B sky130_fd_sc_hd__a221oi_2
XPHY_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _13608_/Q vssd1 vssd1 vccd1 vccd1 _11680_/Y sky130_fd_sc_hd__inv_2
XPHY_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _14295_/Q vssd1 vssd1 vccd1 vccd1 _10631_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _13350_/CLK _13350_/D vssd1 vssd1 vccd1 vccd1 _13350_/Q sky130_fd_sc_hd__dfxtp_1
X_10562_ _14060_/Q vssd1 vssd1 vccd1 vccd1 _10562_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _11271_/Y _14542_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13281_ _14573_/CLK _13281_/D vssd1 vssd1 vccd1 vccd1 _13281_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _13583_/Q vssd1 vssd1 vccd1 vccd1 _10493_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12232_ _12232_/A vssd1 vssd1 vccd1 vccd1 _12232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12163_ vssd1 vssd1 vccd1 vccd1 _12163_/HI _12163_/LO sky130_fd_sc_hd__conb_1
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _14461_/Q vssd1 vssd1 vccd1 vccd1 _11114_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12094_ vssd1 vssd1 vccd1 vccd1 _12094_/HI _12094_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11045_ _13953_/Q vssd1 vssd1 vccd1 vccd1 _11045_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _12578_/X input343/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11947_ _11928_/X _11947_/B _11947_/C _11947_/D vssd1 vssd1 vccd1 vccd1 _11948_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _11876_/Y _10181_/A _11877_/Y _10184_/A vssd1 vssd1 vccd1 vccd1 _11878_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13617_ _14047_/CLK _13617_/D vssd1 vssd1 vccd1 vccd1 _13617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10829_ _14260_/Q vssd1 vssd1 vccd1 vccd1 _10829_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ _14621_/CLK _14597_/D vssd1 vssd1 vccd1 vccd1 _14597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13548_ _14120_/CLK _13548_/D vssd1 vssd1 vccd1 vccd1 _13548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13479_ _14188_/CLK _13479_/D vssd1 vssd1 vccd1 vccd1 _13479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07971_ _14084_/Q _07965_/X _07825_/X _07967_/X _07970_/X vssd1 vssd1 vccd1 vccd1
+ _14084_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09710_ _09707_/X _09709_/X _09707_/X _09709_/X vssd1 vssd1 vccd1 vccd1 _09710_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06922_ _06919_/X _12299_/X _06920_/Y _06921_/X vssd1 vssd1 vccd1 vccd1 _06923_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09641_ _09641_/A vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06853_ _06853_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _06853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ _09570_/X _09569_/X _13266_/Q _09571_/X vssd1 vssd1 vccd1 vccd1 _13234_/D
+ sky130_fd_sc_hd__o22a_1
X_06784_ _08146_/A vssd1 vssd1 vccd1 vccd1 _06784_/X sky130_fd_sc_hd__buf_2
XFILLER_208_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08523_ _08927_/A vssd1 vssd1 vccd1 vccd1 _08523_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08454_ _13837_/Q _08452_/X _08150_/X _08453_/X _08449_/X vssd1 vssd1 vccd1 vccd1
+ _13837_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07405_ _14365_/Q _07307_/A _07083_/X _07309_/A _07397_/X vssd1 vssd1 vccd1 vccd1
+ _14365_/D sky130_fd_sc_hd__o221a_1
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08385_ _13874_/Q _08379_/X _08155_/X _08380_/X _08384_/X vssd1 vssd1 vccd1 vccd1
+ _13874_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07336_ _08123_/A vssd1 vssd1 vccd1 vccd1 _07336_/X sky130_fd_sc_hd__buf_2
XFILLER_104_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07267_ _14427_/Q _07265_/X _06771_/X _07266_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _14427_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09006_ _09040_/A vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07198_ _14464_/Q _07193_/X _06778_/X _07194_/X _07197_/X vssd1 vssd1 vccd1 vccd1
+ _14464_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _13312_/Q vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__inv_2
XFILLER_134_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09839_ _13330_/Q _09837_/Y _09781_/B vssd1 vssd1 vccd1 vccd1 _09839_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _12523_/X _12849_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12850_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11791_/Y _11646_/X _11794_/X _11797_/X _11800_/X vssd1 vssd1 vccd1 vccd1
+ _11823_/C sky130_fd_sc_hd__o2111a_4
XPHY_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _09526_/X _12780_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__mux2_1
XPHY_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14637_/CLK _14520_/D vssd1 vssd1 vccd1 vccd1 _14520_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11732_ _11727_/Y _11679_/X _11728_/Y _11681_/X _11731_/X vssd1 vssd1 vccd1 vccd1
+ _11739_/C sky130_fd_sc_hd__o221a_1
XPHY_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14529_/CLK _14451_/D vssd1 vssd1 vccd1 vccd1 _14451_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11663_/A vssd1 vssd1 vccd1 vccd1 _11663_/X sky130_fd_sc_hd__buf_2
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13402_ _14188_/CLK _13402_/D vssd1 vssd1 vccd1 vccd1 _13402_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10614_ _13866_/Q vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__inv_2
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _14627_/CLK _14382_/D vssd1 vssd1 vccd1 vccd1 _14382_/Q sky130_fd_sc_hd__dfxtp_1
X_11594_ _13646_/Q vssd1 vssd1 vccd1 vccd1 _11594_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13333_ _13352_/CLK _13333_/D vssd1 vssd1 vccd1 vccd1 _13333_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10545_ _14371_/Q vssd1 vssd1 vccd1 vccd1 _10545_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13264_ _14639_/CLK _13264_/D vssd1 vssd1 vccd1 vccd1 _13264_/Q sky130_fd_sc_hd__dfxtp_2
X_10476_ _14487_/Q vssd1 vssd1 vccd1 vccd1 _10476_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12215_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _14071_/CLK _13195_/D vssd1 vssd1 vccd1 vccd1 _13195_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12146_ vssd1 vssd1 vccd1 vccd1 _12146_/HI _12146_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ vssd1 vssd1 vccd1 vccd1 _12077_/HI _12077_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11028_ _13913_/Q vssd1 vssd1 vccd1 vccd1 _11028_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12979_ _12568_/X _12978_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12979_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_16 _11740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_27 _08126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08170_ _13985_/Q _08161_/X _08169_/X _08163_/X _08159_/X vssd1 vssd1 vccd1 vccd1
+ _13985_/D sky130_fd_sc_hd__o221a_1
XANTENNA_38 _06850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _07712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07121_ _14505_/Q _07119_/X _06771_/X _07120_/X _07114_/X vssd1 vssd1 vccd1 vccd1
+ _14505_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07052_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _08007_/A vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__clkbuf_2
XPHY_6908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06905_ _06917_/A _06905_/B vssd1 vssd1 vccd1 vccd1 _14588_/D sky130_fd_sc_hd__nor2_1
X_07885_ _14130_/Q _07882_/X _07809_/X _07884_/X _07872_/X vssd1 vssd1 vccd1 vccd1
+ _14130_/D sky130_fd_sc_hd__o221a_1
X_09624_ _14583_/Q _14565_/Q _06920_/Y _06985_/Y vssd1 vssd1 vccd1 vccd1 _09624_/X
+ sky130_fd_sc_hd__o22a_1
X_06836_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08183_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _09544_/X _09554_/X _13272_/Q _09545_/X vssd1 vssd1 vccd1 vccd1 _13240_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06767_ _06785_/A vssd1 vssd1 vccd1 vccd1 _06767_/X sky130_fd_sc_hd__buf_2
XFILLER_58_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08506_ _13812_/Q _08500_/X _08505_/X _08503_/X _08497_/X vssd1 vssd1 vccd1 vccd1
+ _13812_/D sky130_fd_sc_hd__o221a_1
XFILLER_93_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09486_ _09500_/A vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__clkbuf_2
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06698_ _08922_/A _06697_/X _08922_/A _06697_/X vssd1 vssd1 vccd1 vccd1 _06698_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08437_/X sky130_fd_sc_hd__clkbuf_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08368_ _13884_/Q _08363_/X _08128_/X _08364_/X _08367_/X vssd1 vssd1 vccd1 vccd1
+ _13884_/D sky130_fd_sc_hd__o221a_1
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07319_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07319_/X sky130_fd_sc_hd__buf_2
XFILLER_176_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ _13923_/Q _08293_/X _08128_/X _08294_/X _08297_/X vssd1 vssd1 vccd1 vccd1
+ _13923_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ _14250_/Q vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10261_ _10256_/Y _10150_/X _10257_/Y _10153_/X _10260_/X vssd1 vssd1 vccd1 vccd1
+ _10298_/A sky130_fd_sc_hd__o221a_2
XFILLER_156_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _13896_/Q vssd1 vssd1 vccd1 vccd1 _12000_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _10186_/Y _10188_/X _10189_/Y _10191_/X vssd1 vssd1 vccd1 vccd1 _10192_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13951_ _14107_/CLK _13951_/D vssd1 vssd1 vccd1 vccd1 _13951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12902_ _12536_/X _12901_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13882_ _14110_/CLK _13882_/D vssd1 vssd1 vccd1 vccd1 _13882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12833_ _12519_/X _12832_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12833_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12764_ _09509_/X input354/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12764_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _14006_/Q vssd1 vssd1 vccd1 vccd1 _11715_/Y sky130_fd_sc_hd__inv_2
X_14503_ _14621_/CLK _14503_/D vssd1 vssd1 vccd1 vccd1 _14503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12695_ _09595_/X _12694_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13192_/D sky130_fd_sc_hd__mux2_1
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11646_ _11646_/A vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__buf_2
X_14434_ _14527_/CLK _14434_/D vssd1 vssd1 vccd1 vccd1 _14434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 io_in[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 io_in[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
X_14365_ _14633_/CLK _14365_/D vssd1 vssd1 vccd1 vccd1 _14365_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 io_in[7] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XFILLER_200_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11577_ _14315_/Q vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput47 la_data_in[107] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_1
Xinput58 la_data_in[117] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
X_13316_ _14538_/CLK _13316_/D vssd1 vssd1 vccd1 vccd1 _13316_/Q sky130_fd_sc_hd__dfxtp_1
X_10528_ _13942_/Q vssd1 vssd1 vccd1 vccd1 _10528_/Y sky130_fd_sc_hd__inv_2
Xinput69 la_data_in[127] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14296_ _14305_/CLK _14296_/D vssd1 vssd1 vccd1 vccd1 _14296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13247_ _14538_/CLK _13247_/D vssd1 vssd1 vccd1 vccd1 _13279_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10459_ _10453_/Y _10455_/X _10456_/Y _10458_/X vssd1 vssd1 vccd1 vccd1 _10459_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ _13177_/X _12667_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12129_ vssd1 vssd1 vccd1 vccd1 _12129_/HI _12129_/LO sky130_fd_sc_hd__conb_1
XFILLER_65_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater615 _13114_/S vssd1 vssd1 vccd1 vccd1 _13146_/S sky130_fd_sc_hd__buf_8
XFILLER_61_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater626 _06785_/A vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__buf_6
XFILLER_26_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater637 _13099_/S vssd1 vssd1 vccd1 vccd1 _13147_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater648 _14527_/CLK vssd1 vssd1 vccd1 vccd1 _14637_/CLK sky130_fd_sc_hd__buf_12
XFILLER_61_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater659 _14056_/CLK vssd1 vssd1 vccd1 vccd1 _14169_/CLK sky130_fd_sc_hd__buf_12
XFILLER_113_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07670_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06621_ _06616_/X _06620_/X _06616_/X _06620_/X vssd1 vssd1 vccd1 vccd1 _06621_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ _09352_/A vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06552_ _06554_/A vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09271_ _09271_/A _09271_/B _09271_/C _09271_/D vssd1 vssd1 vccd1 vccd1 _10168_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_179_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08222_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08222_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08153_ _08153_/A vssd1 vssd1 vccd1 vccd1 _08153_/X sky130_fd_sc_hd__buf_4
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07104_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07104_/X sky130_fd_sc_hd__clkbuf_2
X_08084_ _14019_/Q _08078_/X _07790_/X _08079_/X _08083_/X vssd1 vssd1 vccd1 vccd1
+ _14019_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _07061_/A vssd1 vssd1 vccd1 vccd1 _07035_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08986_/X sky130_fd_sc_hd__clkbuf_4
XPHY_7439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07937_ _09535_/A vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__clkbuf_4
XPHY_6738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07868_ _14138_/Q _07863_/X _07867_/X _07864_/X _07865_/X vssd1 vssd1 vccd1 vccd1
+ _14138_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06819_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08171_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09607_ _09607_/A vssd1 vssd1 vccd1 vccd1 _12974_/S sky130_fd_sc_hd__buf_2
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07799_ _14172_/Q _07704_/A _07798_/X _07706_/A _07794_/X vssd1 vssd1 vccd1 vccd1
+ _14172_/D sky130_fd_sc_hd__o221a_1
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ _09530_/X _09537_/X _13279_/Q _09531_/X vssd1 vssd1 vccd1 vccd1 _13247_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _13284_/Q _09464_/X _12279_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _13284_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _13923_/Q vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__inv_2
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12479_/X _06961_/Y _12486_/S vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11431_/A vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _14305_/CLK _14150_/D vssd1 vssd1 vccd1 vccd1 _14150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11362_ _14233_/Q _11170_/X _14428_/Q _11171_/X _11361_/X vssd1 vssd1 vccd1 vccd1
+ _11395_/B sky130_fd_sc_hd__a221oi_2
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _12629_/X _13100_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _13101_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10313_ _14094_/Q vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ _14529_/CLK _14081_/D vssd1 vssd1 vccd1 vccd1 _14081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11293_ _13213_/Q _11249_/X _14036_/Q _11193_/X _11292_/X vssd1 vssd1 vccd1 vccd1
+ _11293_/X sky130_fd_sc_hd__a221o_4
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _12596_/X input350/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__mux2_1
X_10244_ _11691_/A vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ _14209_/Q _10164_/X _14404_/Q _10167_/X _10174_/X vssd1 vssd1 vccd1 vccd1
+ _10255_/B sky130_fd_sc_hd__a221oi_2
XFILLER_26_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13934_ _14169_/CLK _13934_/D vssd1 vssd1 vccd1 vccd1 _13934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _14100_/CLK _13865_/D vssd1 vssd1 vccd1 vccd1 _13865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12816_ _12516_/X input352/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ _14114_/CLK _13796_/D vssd1 vssd1 vccd1 vccd1 _13796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12747_ _09547_/X _12746_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13211_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _09586_/X _12677_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12678_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11629_ _11624_/Y _11455_/X _11625_/Y _11457_/X _11628_/X vssd1 vssd1 vccd1 vccd1
+ _11630_/D sky130_fd_sc_hd__o221a_1
X_14417_ _14470_/CLK _14417_/D vssd1 vssd1 vccd1 vccd1 _14417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14348_ _14495_/CLK _14348_/D vssd1 vssd1 vccd1 vccd1 _14348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14279_ _14637_/CLK _14279_/D vssd1 vssd1 vccd1 vccd1 _14279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08840_ _13649_/Q _08832_/X _08837_/X _08835_/X _08839_/X vssd1 vssd1 vccd1 vccd1
+ _13649_/D sky130_fd_sc_hd__o221a_1
XFILLER_83_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08771_ _13683_/Q _08767_/X _08517_/X _08768_/X _08769_/X vssd1 vssd1 vccd1 vccd1
+ _13683_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07722_ _14203_/Q _07718_/X _07719_/X _07721_/X _07715_/X vssd1 vssd1 vccd1 vccd1
+ _14203_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07653_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06604_ _06600_/Y _08957_/A _08948_/A _06603_/Y vssd1 vssd1 vccd1 vccd1 _06604_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07584_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__buf_4
XFILLER_20_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _13394_/Q _09318_/X _08167_/A _09319_/X _09322_/X vssd1 vssd1 vccd1 vccd1
+ _13394_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ _06535_/A vssd1 vssd1 vccd1 vccd1 _06535_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09254_ _13433_/Q _09249_/X _08962_/X _09250_/X _09252_/X vssd1 vssd1 vccd1 vccd1
+ _13433_/D sky130_fd_sc_hd__o221a_1
XFILLER_72_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08205_ _13974_/Q _08198_/X _08199_/X _08201_/X _08204_/X vssd1 vssd1 vccd1 vccd1
+ _13974_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09185_ _13472_/Q _09179_/X _08962_/X _09180_/X _09182_/X vssd1 vssd1 vccd1 vccd1
+ _13472_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08136_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08067_ _14029_/Q _08061_/X _07852_/X _08062_/X _08066_/X vssd1 vssd1 vccd1 vccd1
+ _14029_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07018_ _07028_/A vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput204 la_oenb[18] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__buf_1
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 la_oenb[28] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_1
XPHY_7236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput226 la_oenb[38] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__buf_1
XPHY_7247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 la_oenb[48] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_1
XPHY_7258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput248 la_oenb[58] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__buf_1
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput259 la_oenb[68] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_hd__buf_1
XFILLER_40_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _11978_/Y _10234_/A _11979_/Y _10237_/A vssd1 vssd1 vccd1 vccd1 _11980_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931_ _10922_/Y _10923_/X _10924_/Y _10925_/X _10930_/X vssd1 vssd1 vccd1 vccd1
+ _10993_/A sky130_fd_sc_hd__o221a_4
XPHY_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13650_ _14139_/CLK _13650_/D vssd1 vssd1 vccd1 vccd1 _13650_/Q sky130_fd_sc_hd__dfxtp_1
X_10862_ _14339_/Q vssd1 vssd1 vccd1 vccd1 _10862_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12601_ _09910_/X _13312_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _14173_/CLK _13581_/D vssd1 vssd1 vccd1 vccd1 _13581_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _14454_/Q vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _13368_/Q _10031_/X _12647_/S vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12463_ _12462_/X _06933_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12463_/X sky130_fd_sc_hd__mux2_2
XFILLER_16_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ _14481_/CLK _14202_/D vssd1 vssd1 vccd1 vccd1 _14202_/Q sky130_fd_sc_hd__dfxtp_1
X_11414_ _11414_/A vssd1 vssd1 vccd1 vccd1 _11414_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12394_ _12393_/X _13207_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14133_ _14173_/CLK _14133_/D vssd1 vssd1 vccd1 vccd1 _14133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11345_ _11343_/Y _11213_/X _11344_/Y _11215_/X vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14064_ _14119_/CLK _14064_/D vssd1 vssd1 vccd1 vccd1 _14064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11276_ _11274_/Y _11165_/X _11275_/Y _11167_/X vssd1 vssd1 vccd1 vccd1 _11276_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_165_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13015_ _12586_/X _13014_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _11679_/A vssd1 vssd1 vccd1 vccd1 _10228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _11639_/A vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10089_ _12510_/S _10089_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__or2_2
XFILLER_43_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13917_ _14146_/CLK _13917_/D vssd1 vssd1 vccd1 vccd1 _13917_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _14094_/CLK _13848_/D vssd1 vssd1 vccd1 vccd1 _13848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _14130_/CLK _13779_/D vssd1 vssd1 vccd1 vccd1 _13779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09941_ _09903_/A _09903_/B _09940_/Y vssd1 vssd1 vccd1 vccd1 _09941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09872_ _13296_/Q vssd1 vssd1 vccd1 vccd1 _09890_/A sky130_fd_sc_hd__inv_2
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08823_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08823_/X sky130_fd_sc_hd__buf_2
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08754_ _13692_/Q _08748_/X _08492_/X _08750_/X _08751_/X vssd1 vssd1 vccd1 vccd1
+ _13692_/D sky130_fd_sc_hd__o221a_1
XPHY_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07705_ _07785_/A vssd1 vssd1 vccd1 vccd1 _07706_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08685_ _13729_/Q _08677_/X _08496_/X _08679_/X _08684_/X vssd1 vssd1 vccd1 vccd1
+ _13729_/D sky130_fd_sc_hd__o221a_1
XPHY_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07636_/A vssd1 vssd1 vccd1 vccd1 _07636_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07567_ _14284_/Q _07561_/X _07313_/X _07563_/X _07566_/X vssd1 vssd1 vccd1 vccd1
+ _14284_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09306_ _09306_/A vssd1 vssd1 vccd1 vccd1 _09306_/X sky130_fd_sc_hd__clkbuf_2
X_06518_ _06853_/A _09732_/A vssd1 vssd1 vccd1 vccd1 _08813_/A sky130_fd_sc_hd__or2_4
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _07541_/A vssd1 vssd1 vccd1 vccd1 _07532_/A sky130_fd_sc_hd__buf_4
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _13444_/Q _09233_/X _08933_/X _09234_/X _09236_/X vssd1 vssd1 vccd1 vccd1
+ _13444_/D sky130_fd_sc_hd__o221a_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09168_ _13482_/Q _09163_/X _08935_/X _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1
+ _13482_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08119_ _08119_/A vssd1 vssd1 vccd1 vccd1 _08119_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09099_ _13521_/Q _09095_/X _08935_/X _09096_/X _09093_/X vssd1 vssd1 vccd1 vccd1
+ _13521_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _11128_/Y _10942_/X _11129_/Y _10944_/X vssd1 vssd1 vccd1 vccd1 _11130_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11061_ _14382_/Q vssd1 vssd1 vccd1 vccd1 _11061_/Y sky130_fd_sc_hd__inv_2
XPHY_7000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10012_ _13376_/Q _10011_/B _10013_/A vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__o21a_1
XPHY_7033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _11961_/Y _10188_/A _11962_/Y _10191_/A vssd1 vssd1 vccd1 vccd1 _11963_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _14178_/CLK _13702_/D vssd1 vssd1 vccd1 vccd1 _13702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10914_ _13911_/Q vssd1 vssd1 vccd1 vccd1 _10914_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11894_ _14322_/Q vssd1 vssd1 vccd1 vccd1 _11894_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13633_ _14071_/CLK _13633_/D vssd1 vssd1 vccd1 vccd1 _13633_/Q sky130_fd_sc_hd__dfxtp_1
X_10845_ _10840_/Y _10687_/X _10841_/Y _10689_/X _10844_/X vssd1 vssd1 vccd1 vccd1
+ _10880_/A sky130_fd_sc_hd__o221a_2
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13564_ _14120_/CLK _13564_/D vssd1 vssd1 vccd1 vccd1 _13564_/Q sky130_fd_sc_hd__dfxtp_1
X_10776_ _13550_/Q _10720_/X _13791_/Q _10721_/X vssd1 vssd1 vccd1 vccd1 _10776_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12515_ _13354_/Q _10052_/Y _12610_/S vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__mux2_1
X_13495_ _14173_/CLK _13495_/D vssd1 vssd1 vccd1 vccd1 _13495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12446_ _12509_/X _06915_/Y _12446_/S vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput508 _12102_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__clkbuf_2
X_12377_ _13212_/Q _06596_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput519 _12103_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14116_ _14119_/CLK _14116_/D vssd1 vssd1 vccd1 vccd1 _14116_/Q sky130_fd_sc_hd__dfxtp_1
X_11328_ _11326_/Y _11183_/X _11327_/Y _11185_/X vssd1 vssd1 vccd1 vccd1 _11328_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14047_ _14047_/CLK _14047_/D vssd1 vssd1 vccd1 vccd1 _14047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11259_ _13599_/Q vssd1 vssd1 vccd1 vccd1 _11259_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08470_ _13827_/Q _08468_/X _08175_/X _08469_/X _08465_/X vssd1 vssd1 vccd1 vccd1
+ _13827_/D sky130_fd_sc_hd__o221a_1
XFILLER_93_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07421_ _07467_/A vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ _08140_/A vssd1 vssd1 vccd1 vccd1 _07352_/X sky130_fd_sc_hd__buf_2
XFILLER_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _09039_/A vssd1 vssd1 vccd1 vccd1 _09022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09924_ _13316_/Q _09920_/Y _09926_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09855_ _13325_/Q _09853_/Y _09776_/B vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08806_ _13661_/Q _08800_/X _08572_/X _08801_/X _08802_/X vssd1 vssd1 vccd1 vccd1
+ _13661_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09786_ _09786_/A _09820_/A vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__or2_2
X_06998_ _07004_/A _06998_/B vssd1 vssd1 vccd1 vccd1 _14562_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08737_ _08777_/A vssd1 vssd1 vccd1 vccd1 _08737_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 _10211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _10583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_128 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _13737_/Q _08662_/X _08494_/X _08663_/X _08665_/X vssd1 vssd1 vccd1 vccd1
+ _13737_/D sky130_fd_sc_hd__o221a_1
XPHY_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _11487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07619_ _14253_/Q _07613_/X _07394_/X _07614_/X _07617_/X vssd1 vssd1 vccd1 vccd1
+ _14253_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08599_ _08635_/A vssd1 vssd1 vccd1 vccd1 _08599_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10630_ _10625_/Y _10478_/X _10626_/Y _10481_/X _10629_/X vssd1 vssd1 vccd1 vccd1
+ _10643_/B sky130_fd_sc_hd__o221a_2
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10561_ _10561_/A _10561_/B _10561_/C _10561_/D vssd1 vssd1 vccd1 vccd1 _10561_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_17_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12300_ _11313_/Y _14543_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _14538_/CLK _13280_/D vssd1 vssd1 vccd1 vccd1 _13280_/Q sky130_fd_sc_hd__dfxtp_4
X_10492_ _11445_/A vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ vssd1 vssd1 vccd1 vccd1 _12162_/HI _12162_/LO sky130_fd_sc_hd__conb_1
XFILLER_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11113_ _13479_/Q vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12093_ vssd1 vssd1 vccd1 vccd1 _12093_/HI _12093_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11044_ _14226_/Q _10933_/X _14421_/Q _10935_/X _11043_/X vssd1 vssd1 vccd1 vccd1
+ _11077_/B sky130_fd_sc_hd__a221oi_2
XFILLER_150_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12995_ _12576_/X _12994_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _11941_/Y _10242_/A _11942_/Y _10245_/A _11945_/X vssd1 vssd1 vccd1 vccd1
+ _11947_/D sky130_fd_sc_hd__o221a_1
XPHY_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11877_ _13893_/Q vssd1 vssd1 vccd1 vccd1 _11877_/Y sky130_fd_sc_hd__inv_2
XPHY_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ _14173_/CLK _13616_/D vssd1 vssd1 vccd1 vccd1 _13616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ _14182_/Q vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14596_ _14621_/CLK _14596_/D vssd1 vssd1 vccd1 vccd1 _14596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13547_ _14121_/CLK _13547_/D vssd1 vssd1 vccd1 vccd1 _13547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10759_ _13628_/Q vssd1 vssd1 vccd1 vccd1 _10759_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13478_ _14188_/CLK _13478_/D vssd1 vssd1 vccd1 vccd1 _13478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12429_ _12428_/X _06893_/X _12603_/S vssd1 vssd1 vccd1 vccd1 _12429_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _07978_/A vssd1 vssd1 vccd1 vccd1 _07970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06921_ _06958_/A vssd1 vssd1 vccd1 vccd1 _06921_/X sky130_fd_sc_hd__buf_1
XFILLER_136_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06852_ _14599_/Q _06530_/A _06716_/X _08268_/A _06838_/X vssd1 vssd1 vccd1 vccd1
+ _14599_/D sky130_fd_sc_hd__o221a_1
X_09640_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06783_ _08942_/A vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08522_ _13805_/Q _08513_/X _08521_/X _08515_/X _08511_/X vssd1 vssd1 vccd1 vccd1
+ _13805_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08453_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07404_ _14366_/Q _07307_/A _07403_/X _07309_/A _07397_/X vssd1 vssd1 vccd1 vccd1
+ _14366_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08384_ _08421_/A vssd1 vssd1 vccd1 vccd1 _08384_/X sky130_fd_sc_hd__buf_2
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07335_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07335_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07266_ _07283_/A vssd1 vssd1 vccd1 vccd1 _07266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09005_ _09049_/A vssd1 vssd1 vccd1 vccd1 _09040_/A sky130_fd_sc_hd__buf_2
XFILLER_121_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07197_ _07213_/A vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__buf_2
XFILLER_195_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _09905_/A _09905_/B _09906_/Y vssd1 vssd1 vccd1 vccd1 _09907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09838_ _09779_/A _09779_/B _09837_/Y vssd1 vssd1 vccd1 vccd1 _09838_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _13319_/Q vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__inv_2
XFILLER_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11798_/Y _11658_/X _11799_/Y _11660_/X vssd1 vssd1 vccd1 vccd1 _11800_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _09526_/X input349/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12780_/X sky130_fd_sc_hd__mux2_1
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11729_/Y _11683_/X _11730_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11731_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14529_/CLK _14450_/D vssd1 vssd1 vccd1 vccd1 _14450_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11662_ _11645_/Y _11646_/X _11651_/X _11656_/X _11661_/X vssd1 vssd1 vccd1 vccd1
+ _11699_/C sky130_fd_sc_hd__o2111a_4
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _14188_/CLK _13401_/D vssd1 vssd1 vccd1 vccd1 _13401_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10613_ _13749_/Q vssd1 vssd1 vccd1 vccd1 _10613_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _13685_/Q vssd1 vssd1 vccd1 vccd1 _11593_/Y sky130_fd_sc_hd__inv_2
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _14627_/CLK _14381_/D vssd1 vssd1 vccd1 vccd1 _14381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10544_ _14605_/Q vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__inv_2
X_13332_ _13877_/CLK _13332_/D vssd1 vssd1 vccd1 vccd1 _13332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ _13196_/Q _10276_/X _14019_/Q _10469_/X _10474_/X vssd1 vssd1 vccd1 vccd1
+ _10475_/X sky130_fd_sc_hd__a221o_4
XFILLER_13_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13263_ _14639_/CLK _13263_/D vssd1 vssd1 vccd1 vccd1 _13263_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12214_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13194_ _14114_/CLK _13194_/D vssd1 vssd1 vccd1 vccd1 _13194_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12145_ vssd1 vssd1 vccd1 vccd1 _12145_/HI _12145_/LO sky130_fd_sc_hd__conb_1
XFILLER_151_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12076_ vssd1 vssd1 vccd1 vccd1 _12076_/HI _12076_/LO sky130_fd_sc_hd__conb_1
XFILLER_133_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11027_ _11022_/Y _10973_/X _11023_/Y _10975_/X _11026_/X vssd1 vssd1 vccd1 vccd1
+ _11034_/C sky130_fd_sc_hd__o221a_1
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ _12977_/X _12568_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11929_ _14518_/Q vssd1 vssd1 vccd1 vccd1 _11929_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_17 _11782_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_28 _08137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_39 _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14579_ _14621_/CLK _14579_/D vssd1 vssd1 vccd1 vccd1 _14579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07051_ _14540_/Q _07044_/X _06784_/X _07045_/X _07046_/X vssd1 vssd1 vccd1 vccd1
+ _14540_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07953_ _08008_/A vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__inv_2
XFILLER_9_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06904_ _06901_/X _12294_/X _06902_/Y _06903_/X vssd1 vssd1 vccd1 vccd1 _06905_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_07884_ _07884_/A vssd1 vssd1 vccd1 vccd1 _07884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09623_ _06943_/X _14562_/Q _14577_/Q _06996_/Y vssd1 vssd1 vccd1 vccd1 _09623_/X
+ sky130_fd_sc_hd__o22a_1
X_06835_ _14604_/Q _06823_/X _06834_/X _06532_/A _06821_/X vssd1 vssd1 vccd1 vccd1
+ _14604_/D sky130_fd_sc_hd__o221a_1
XFILLER_77_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06766_ _08132_/A vssd1 vssd1 vccd1 vccd1 _06766_/X sky130_fd_sc_hd__buf_2
X_09554_ _09560_/A _12391_/X vssd1 vssd1 vccd1 vccd1 _09554_/X sky130_fd_sc_hd__and2_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08505_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09485_ _13272_/Q _09479_/X _12267_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _13272_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06697_ _06600_/Y _06656_/Y _08948_/A _08950_/A vssd1 vssd1 vccd1 vccd1 _06697_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08436_ _08460_/A vssd1 vssd1 vccd1 vccd1 _08436_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08367_/X sky130_fd_sc_hd__buf_2
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07318_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__buf_2
X_08298_ _13924_/Q _08293_/X _08126_/X _08294_/X _08297_/X vssd1 vssd1 vccd1 vccd1
+ _13924_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07249_ _07291_/A vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__buf_4
XFILLER_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _10258_/Y _10156_/X _10259_/Y _10159_/X vssd1 vssd1 vccd1 vccd1 _10260_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10191_ _10191_/A vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _14107_/CLK _13950_/D vssd1 vssd1 vccd1 vccd1 _13950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12901_ _12536_/X _12900_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13881_ _13996_/CLK _13881_/D vssd1 vssd1 vccd1 vccd1 _13881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12832_ _12519_/X input335/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12763_ _09556_/X _12762_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13207_/D sky130_fd_sc_hd__mux2_1
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14502_ _14621_/CLK _14502_/D vssd1 vssd1 vccd1 vccd1 _14502_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11714_ _11712_/Y _11653_/X _11713_/Y _11655_/X vssd1 vssd1 vccd1 vccd1 _11714_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _09595_/X _12693_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__mux2_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14433_ _14527_/CLK _14433_/D vssd1 vssd1 vccd1 vccd1 _14433_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11645_ _13966_/Q vssd1 vssd1 vccd1 vccd1 _11645_/Y sky130_fd_sc_hd__inv_2
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 io_in[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
XFILLER_204_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14364_ _14637_/CLK _14364_/D vssd1 vssd1 vccd1 vccd1 _14364_/Q sky130_fd_sc_hd__dfxtp_1
Xinput26 io_in[32] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XFILLER_141_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11576_ _11571_/Y _11435_/X _11572_/Y _11437_/X _11575_/X vssd1 vssd1 vccd1 vccd1
+ _11589_/B sky130_fd_sc_hd__o221a_2
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 io_in[8] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_1
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 la_data_in[108] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_1
Xinput59 la_data_in[118] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
X_13315_ _14538_/CLK _13315_/D vssd1 vssd1 vccd1 vccd1 _13315_/Q sky130_fd_sc_hd__dfxtp_1
X_10527_ _14215_/Q _10437_/X _14410_/Q _10438_/X _10526_/X vssd1 vssd1 vccd1 vccd1
+ _10561_/B sky130_fd_sc_hd__a221oi_2
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14295_ _14529_/CLK _14295_/D vssd1 vssd1 vccd1 vccd1 _14295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10458_ _11421_/A vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13246_ _14538_/CLK _13246_/D vssd1 vssd1 vccd1 vccd1 _13278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10389_ _14213_/Q _10164_/X _14408_/Q _10167_/X _10388_/X vssd1 vssd1 vccd1 vccd1
+ _10422_/B sky130_fd_sc_hd__a221oi_2
X_13177_ _12667_/X _13176_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12128_ vssd1 vssd1 vccd1 vccd1 _12128_/HI _12128_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12059_ _09788_/A _12057_/X _09900_/A _12058_/X vssd1 vssd1 vccd1 vccd1 _12059_/Y
+ sky130_fd_sc_hd__o22ai_1
Xrepeater616 _13110_/S vssd1 vssd1 vccd1 vccd1 _13114_/S sky130_fd_sc_hd__buf_6
Xrepeater627 _09457_/A vssd1 vssd1 vccd1 vccd1 _06723_/C1 sky130_fd_sc_hd__buf_4
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater638 _14595_/CLK vssd1 vssd1 vccd1 vccd1 _14621_/CLK sky130_fd_sc_hd__buf_12
Xrepeater649 _14527_/CLK vssd1 vssd1 vccd1 vccd1 _14633_/CLK sky130_fd_sc_hd__buf_12
XFILLER_42_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06620_ _06589_/Y _06619_/X _06589_/Y _06619_/X vssd1 vssd1 vccd1 vccd1 _06620_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06551_ _06553_/A vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09270_ _13422_/Q _09205_/A _09060_/X _09207_/A _09267_/X vssd1 vssd1 vccd1 vccd1
+ _13422_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08221_ _08246_/A vssd1 vssd1 vccd1 vccd1 _08221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08152_ _13993_/Q _08149_/X _08150_/X _08151_/X _08147_/X vssd1 vssd1 vccd1 vccd1
+ _13993_/D sky130_fd_sc_hd__o221a_1
XFILLER_72_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07103_ _07145_/A vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__buf_4
XFILLER_200_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08083_ _08120_/A vssd1 vssd1 vccd1 vccd1 _08083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07034_ _14550_/Q _07025_/X _06748_/X _07027_/X _07028_/X vssd1 vssd1 vccd1 vccd1
+ _14550_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ _08985_/A vssd1 vssd1 vccd1 vccd1 _08985_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _14100_/Q _07934_/X _07784_/X _07935_/X _07929_/X vssd1 vssd1 vccd1 vccd1
+ _14100_/D sky130_fd_sc_hd__o221a_1
XPHY_6728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07867_ _08259_/A vssd1 vssd1 vccd1 vccd1 _07867_/X sky130_fd_sc_hd__buf_4
XFILLER_25_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _12035_/A vssd1 vssd1 vccd1 vccd1 _13110_/S sky130_fd_sc_hd__clkbuf_2
X_06818_ _14609_/Q _06805_/X _06817_/X _06811_/X _06803_/X vssd1 vssd1 vccd1 vccd1
+ _14609_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07798_ _08188_/A vssd1 vssd1 vccd1 vccd1 _07798_/X sky130_fd_sc_hd__buf_4
XFILLER_77_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09537_ _09547_/A _12418_/X vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__and2_1
X_06749_ _06785_/A vssd1 vssd1 vccd1 vccd1 _06749_/X sky130_fd_sc_hd__clkbuf_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _13285_/Q _09464_/X _12280_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _13285_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08419_ _13856_/Q _08415_/X _08099_/X _08417_/X _08406_/X vssd1 vssd1 vccd1 vccd1
+ _13856_/D sky130_fd_sc_hd__o221a_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09399_ _09401_/A _13147_/X vssd1 vssd1 vccd1 vccd1 _13335_/D sky130_fd_sc_hd__and2_1
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11430_ _11430_/A vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11361_ _13407_/Q _11278_/X _13719_/Q _11172_/X vssd1 vssd1 vccd1 vccd1 _11361_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10312_ _13821_/Q vssd1 vssd1 vccd1 vccd1 _10312_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ _12629_/X input332/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ _14529_/CLK _14080_/D vssd1 vssd1 vccd1 vccd1 _14080_/Q sky130_fd_sc_hd__dfxtp_1
X_11292_ _13561_/Q _11194_/X _13802_/Q _11195_/X vssd1 vssd1 vccd1 vccd1 _11292_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10243_ _14131_/Q vssd1 vssd1 vccd1 vccd1 _10243_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _12594_/X _13030_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10174_ _13383_/Q _11747_/A _13695_/Q _10173_/X vssd1 vssd1 vccd1 vccd1 _10174_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13933_ _14169_/CLK _13933_/D vssd1 vssd1 vccd1 vccd1 _13933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13864_ _14100_/CLK _13864_/D vssd1 vssd1 vccd1 vccd1 _13864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _12515_/X _12814_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13795_ _14114_/CLK _13795_/D vssd1 vssd1 vccd1 vccd1 _13795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ _09547_/X _12745_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _09586_/X _12676_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__mux2_1
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14416_ _14470_/CLK _14416_/D vssd1 vssd1 vccd1 vccd1 _14416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11628_ _11626_/Y _11459_/X _11627_/Y _11461_/X vssd1 vssd1 vccd1 vccd1 _11628_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14347_ _14495_/CLK _14347_/D vssd1 vssd1 vccd1 vccd1 _14347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11559_ _13769_/Q vssd1 vssd1 vccd1 vccd1 _11559_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14278_ _14637_/CLK _14278_/D vssd1 vssd1 vccd1 vccd1 _14278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _13352_/CLK _13229_/D vssd1 vssd1 vccd1 vccd1 _13261_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08770_ _13684_/Q _08767_/X _08514_/X _08768_/X _08769_/X vssd1 vssd1 vccd1 vccd1
+ _13684_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07721_ _07772_/A vssd1 vssd1 vccd1 vccd1 _07721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07652_ _14238_/Q _07644_/X _07332_/X _07646_/X _07650_/X vssd1 vssd1 vccd1 vccd1
+ _14238_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06603_ _06603_/A vssd1 vssd1 vccd1 vccd1 _06603_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07583_ _14275_/Q _07580_/X _07339_/X _07581_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _14275_/D sky130_fd_sc_hd__o221a_1
XFILLER_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09322_ _09519_/A vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06534_ _06536_/A vssd1 vssd1 vccd1 vccd1 _08837_/A sky130_fd_sc_hd__buf_4
XFILLER_181_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09253_ _13434_/Q _09249_/X _08960_/X _09250_/X _09252_/X vssd1 vssd1 vccd1 vccd1
+ _13434_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09184_ _13473_/Q _09179_/X _08960_/X _09180_/X _09182_/X vssd1 vssd1 vccd1 vccd1
+ _13473_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08135_ _13999_/Q _08122_/X _08132_/X _08124_/X _08134_/X vssd1 vssd1 vccd1 vccd1
+ _13999_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08066_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07017_ _07017_/A vssd1 vssd1 vccd1 vccd1 _07017_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput205 la_oenb[19] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__buf_1
XFILLER_66_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 la_oenb[29] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_1
XPHY_7237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput227 la_oenb[39] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_1
XFILLER_83_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 la_oenb[49] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_1
XPHY_7259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _13587_/Q _08956_/X _08967_/X _08958_/X _08963_/X vssd1 vssd1 vccd1 vccd1
+ _13587_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 la_oenb[59] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__buf_1
XFILLER_25_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ _07927_/A vssd1 vssd1 vccd1 vccd1 _07919_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ _13615_/Q _08894_/X _08822_/X _08897_/X _08886_/X vssd1 vssd1 vccd1 vccd1
+ _13615_/D sky130_fd_sc_hd__o221a_1
XPHY_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10930_ _10926_/Y _10927_/X _10928_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _10930_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10861_ _14495_/Q vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _13313_/Q _12599_/X _12667_/S vssd1 vssd1 vccd1 vccd1 _12600_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13580_ _14173_/CLK _13580_/D vssd1 vssd1 vccd1 vccd1 _13580_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10792_ _13472_/Q vssd1 vssd1 vccd1 vccd1 _10792_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _13369_/Q _10032_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12531_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12462_ _12461_/X _06933_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12462_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ _14481_/CLK _14201_/D vssd1 vssd1 vccd1 vccd1 _14201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11413_ _13766_/Q vssd1 vssd1 vccd1 vccd1 _11413_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12393_ _13207_/Q _12392_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12393_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14173_/CLK _14132_/D vssd1 vssd1 vccd1 vccd1 _14132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11344_ _14271_/Q vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14063_ _14143_/CLK _14063_/D vssd1 vssd1 vccd1 vccd1 _14063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11275_ _13639_/Q vssd1 vssd1 vccd1 vccd1 _11275_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ _13013_/X _12586_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _13014_/X sky130_fd_sc_hd__mux2_1
X_10226_ _14287_/Q vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _13617_/Q vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10088_ _10094_/A _12487_/X vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__nor2_8
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _14146_/CLK _13916_/D vssd1 vssd1 vccd1 vccd1 _13916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13847_ _14094_/CLK _13847_/D vssd1 vssd1 vccd1 vccd1 _13847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ _14130_/CLK _13778_/D vssd1 vssd1 vccd1 vccd1 _13778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12729_ _09578_/X _12728_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _09940_/A vssd1 vssd1 vccd1 vccd1 _09940_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09871_ _13297_/Q vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__inv_2
XFILLER_119_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08822_ _08822_/A vssd1 vssd1 vccd1 vccd1 _08822_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_140_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08753_ _13693_/Q _08748_/X _08490_/X _08750_/X _08751_/X vssd1 vssd1 vccd1 vccd1
+ _13693_/D sky130_fd_sc_hd__o221a_1
XPHY_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07704_ _07704_/A vssd1 vssd1 vccd1 vccd1 _07704_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08684_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08684_/X sky130_fd_sc_hd__buf_2
XPHY_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07635_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07636_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07566_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07566_/X sky130_fd_sc_hd__buf_2
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09305_ _13405_/Q _09302_/X _08140_/A _09303_/X _09298_/X vssd1 vssd1 vccd1 vccd1
+ _13405_/D sky130_fd_sc_hd__o221a_1
X_06517_ _12667_/S vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__buf_6
X_07497_ _14321_/Q _07488_/X _07317_/X _07490_/X _07493_/X vssd1 vssd1 vccd1 vccd1
+ _14321_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09236_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09236_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_210_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09167_ _13483_/Q _09163_/X _08933_/X _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1
+ _13483_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08118_ _14005_/Q _08109_/X _08117_/X _08112_/X _08106_/X vssd1 vssd1 vccd1 vccd1
+ _14005_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09098_ _13522_/Q _09095_/X _08933_/X _09096_/X _09093_/X vssd1 vssd1 vccd1 vccd1
+ _13522_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08049_ _14040_/Q _08045_/X _07738_/X _08046_/X _08042_/X vssd1 vssd1 vccd1 vccd1
+ _14040_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11060_ _14616_/Q vssd1 vssd1 vccd1 vccd1 _11060_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10011_ _13376_/Q _10011_/B vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__nand2_1
XPHY_7023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _14129_/Q vssd1 vssd1 vccd1 vccd1 _11962_/Y sky130_fd_sc_hd__inv_2
XPHY_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13701_ _14178_/CLK _13701_/D vssd1 vssd1 vccd1 vccd1 _13701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ _10908_/Y _10735_/X _10909_/Y _10737_/X _10912_/X vssd1 vssd1 vccd1 vccd1
+ _10920_/C sky130_fd_sc_hd__o221a_1
XPHY_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _11888_/Y _10214_/A _11889_/Y _10217_/A _11892_/X vssd1 vssd1 vccd1 vccd1
+ _11906_/B sky130_fd_sc_hd__o221a_2
XPHY_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13632_ _14071_/CLK _13632_/D vssd1 vssd1 vccd1 vccd1 _13632_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10842_/Y _10691_/X _10843_/Y _10693_/X vssd1 vssd1 vccd1 vccd1 _10844_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ _14120_/CLK _13563_/D vssd1 vssd1 vccd1 vccd1 _13563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10775_ _11013_/A vssd1 vssd1 vccd1 vccd1 _10775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12514_ _13355_/Q _10053_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12514_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13494_ _14481_/CLK _13494_/D vssd1 vssd1 vccd1 vccd1 _13494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12445_ _12444_/X _06912_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12445_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput509 _12139_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__clkbuf_2
X_12376_ _12375_/X _13213_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14115_ _14120_/CLK _14115_/D vssd1 vssd1 vccd1 vccd1 _14115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11327_ _14115_/Q vssd1 vssd1 vccd1 vccd1 _11327_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _14047_/CLK _14046_/D vssd1 vssd1 vccd1 vccd1 _14046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11258_ _14308_/Q vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10209_ _10209_/A vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11189_ _13520_/Q vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07420_ _14360_/Q _07411_/X _07317_/X _07414_/X _07415_/X vssd1 vssd1 vccd1 vccd1
+ _14360_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07351_ _14388_/Q _07348_/X _07349_/X _07350_/X _07346_/X vssd1 vssd1 vccd1 vccd1
+ _14388_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07282_ _07282_/A vssd1 vssd1 vccd1 vccd1 _07282_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09021_ _13563_/Q _09014_/X _08927_/X _09015_/X _09019_/X vssd1 vssd1 vccd1 vccd1
+ _13563_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__or2_1
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09854_ _09774_/A _09774_/B _09853_/Y vssd1 vssd1 vccd1 vccd1 _09854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08805_ _13662_/Q _08800_/X _08570_/X _08801_/X _08802_/X vssd1 vssd1 vccd1 vccd1
+ _13662_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09785_ _09785_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__or2_1
X_06997_ _06857_/A _12320_/X _06996_/Y _06861_/A vssd1 vssd1 vccd1 vccd1 _06998_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08736_ _08879_/A vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__buf_4
XFILLER_6_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_107 _10278_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _10723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _13738_/Q _08662_/X _08492_/X _08663_/X _08665_/X vssd1 vssd1 vccd1 vccd1
+ _13738_/D sky130_fd_sc_hd__o221a_1
XPHY_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _11251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07618_ _14254_/Q _07613_/X _07392_/X _07614_/X _07617_/X vssd1 vssd1 vccd1 vccd1
+ _14254_/D sky130_fd_sc_hd__o221a_1
XPHY_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08598_ _08643_/A vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__clkbuf_4
XPHY_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07549_ _14290_/Q _07488_/A _07399_/X _07490_/A _07544_/X vssd1 vssd1 vccd1 vccd1
+ _14290_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10541_/X _10560_/B _10560_/C _10560_/D vssd1 vssd1 vccd1 vccd1 _10561_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_122_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09219_ _09219_/A vssd1 vssd1 vccd1 vccd1 _09219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _11679_/A vssd1 vssd1 vccd1 vccd1 _11445_/A sky130_fd_sc_hd__buf_4
XFILLER_194_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12230_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12161_ vssd1 vssd1 vccd1 vccd1 _12161_/HI _12161_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11112_ _14149_/Q vssd1 vssd1 vccd1 vccd1 _11112_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12092_ vssd1 vssd1 vccd1 vccd1 _12092_/HI _12092_/LO sky130_fd_sc_hd__conb_1
XFILLER_46_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11043_ _13400_/Q _11042_/X _13712_/Q _10936_/X vssd1 vssd1 vccd1 vccd1 _11043_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _12993_/X _12576_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11945_ _11943_/Y _10248_/A _11944_/Y _10251_/A vssd1 vssd1 vccd1 vccd1 _11945_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _13776_/Q vssd1 vssd1 vccd1 vccd1 _11876_/Y sky130_fd_sc_hd__inv_2
XPHY_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13615_ _14173_/CLK _13615_/D vssd1 vssd1 vccd1 vccd1 _13615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10827_ _13590_/Q vssd1 vssd1 vccd1 vccd1 _10827_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14595_ _14595_/CLK _14595_/D vssd1 vssd1 vccd1 vccd1 _14595_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13546_ _14121_/CLK _13546_/D vssd1 vssd1 vccd1 vccd1 _13546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10758_ _13667_/Q vssd1 vssd1 vccd1 vccd1 _10758_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13477_ _14188_/CLK _13477_/D vssd1 vssd1 vccd1 vccd1 _13477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10689_ _11399_/A vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12428_ _12509_/X _06893_/X _12428_/S vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ _13202_/Q input99/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06920_ _14583_/Q vssd1 vssd1 vccd1 vccd1 _06920_/Y sky130_fd_sc_hd__inv_2
X_14029_ _14119_/CLK _14029_/D vssd1 vssd1 vccd1 vccd1 _14029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06851_ _09060_/A vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__buf_4
XFILLER_68_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _09583_/A vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__buf_1
X_06782_ _14619_/Q _06769_/X _06781_/X _06772_/X _06767_/X vssd1 vssd1 vccd1 vccd1
+ _14619_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08521_ _08925_/A vssd1 vssd1 vccd1 vccd1 _08521_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08452_ _08460_/A vssd1 vssd1 vccd1 vccd1 _08452_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07403_ _08190_/A vssd1 vssd1 vccd1 vccd1 _07403_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_166_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08383_ _08383_/A vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07334_ _14394_/Q _07322_/X _07332_/X _07325_/X _07333_/X vssd1 vssd1 vccd1 vccd1
+ _14394_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07265_ _07282_/A vssd1 vssd1 vccd1 vccd1 _07265_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09004_ _09039_/A vssd1 vssd1 vccd1 vccd1 _09004_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07196_ _14465_/Q _07193_/X _06775_/X _07194_/X _07189_/X vssd1 vssd1 vccd1 vccd1
+ _14465_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09906_ _09909_/B vssd1 vssd1 vccd1 vccd1 _09906_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _09837_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _13320_/Q vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__inv_2
XPHY_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _13710_/Q _08714_/X _08632_/X _08715_/X _08712_/X vssd1 vssd1 vccd1 vccd1
+ _13710_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09699_ _14568_/Q _06979_/Y _06975_/Y _14567_/Q vssd1 vssd1 vccd1 vccd1 _09699_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _14279_/Q vssd1 vssd1 vccd1 vccd1 _11730_/Y sky130_fd_sc_hd__inv_2
XPHY_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11661_ _11657_/Y _11658_/X _11659_/Y _11660_/X vssd1 vssd1 vccd1 vccd1 _11661_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _14188_/CLK _13400_/D vssd1 vssd1 vccd1 vccd1 _13400_/Q sky130_fd_sc_hd__dfxtp_1
X_10612_ _13944_/Q vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__inv_2
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _14627_/CLK _14380_/D vssd1 vssd1 vccd1 vccd1 _14380_/Q sky130_fd_sc_hd__dfxtp_1
X_11592_ _13451_/Q vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13331_ _14639_/CLK _13331_/D vssd1 vssd1 vccd1 vccd1 _13331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ _14332_/Q vssd1 vssd1 vccd1 vccd1 _10543_/Y sky130_fd_sc_hd__inv_2
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ _14639_/CLK _13262_/D vssd1 vssd1 vccd1 vccd1 _13262_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _13544_/Q _10471_/X _13785_/Q _10473_/X vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12213_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _14071_/CLK _13193_/D vssd1 vssd1 vccd1 vccd1 _13193_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12144_ vssd1 vssd1 vccd1 vccd1 _12144_/HI _12144_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12075_ vssd1 vssd1 vccd1 vccd1 _12075_/HI _12075_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ _11024_/Y _10977_/X _11025_/Y _10979_/X vssd1 vssd1 vccd1 vccd1 _11026_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12977_ _12568_/X _12976_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11928_ _13731_/Q _10173_/A _14050_/Q _10203_/A _11927_/X vssd1 vssd1 vccd1 vccd1
+ _11928_/X sky130_fd_sc_hd__a221o_2
XFILLER_59_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11859_ _13931_/Q vssd1 vssd1 vccd1 vccd1 _11859_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_18 _11823_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14578_ _14621_/CLK _14578_/D vssd1 vssd1 vccd1 vccd1 _14578_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_29 _08146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13529_ _14121_/CLK _13529_/D vssd1 vssd1 vccd1 vccd1 _13529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07050_ _14541_/Q _07044_/X _06781_/X _07045_/X _07046_/X vssd1 vssd1 vccd1 vccd1
+ _14541_/D sky130_fd_sc_hd__o221a_1
XFILLER_12_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07952_ _07952_/A _11633_/A vssd1 vssd1 vccd1 vccd1 _08008_/A sky130_fd_sc_hd__or2_2
XFILLER_155_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06903_ _06958_/A vssd1 vssd1 vccd1 vccd1 _06903_/X sky130_fd_sc_hd__buf_1
XFILLER_151_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07883_ _07935_/A vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__buf_2
XFILLER_25_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09622_ _06993_/Y _09621_/X _06993_/Y _09621_/X vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06834_ _08181_/A vssd1 vssd1 vccd1 vccd1 _06834_/X sky130_fd_sc_hd__buf_2
XFILLER_99_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09544_/X _09552_/X _13273_/Q _09545_/X vssd1 vssd1 vccd1 vccd1 _13241_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06765_ _08927_/A vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__buf_4
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08504_ _13813_/Q _08500_/X _08501_/X _08503_/X _08497_/X vssd1 vssd1 vccd1 vccd1
+ _13813_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09484_ _13273_/Q _09479_/X _12268_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _13273_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06696_ _06696_/A vssd1 vssd1 vccd1 vccd1 _08922_/A sky130_fd_sc_hd__buf_2
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08435_ _13848_/Q _08425_/X _08119_/X _08427_/X _08433_/X vssd1 vssd1 vccd1 vccd1
+ _13848_/D sky130_fd_sc_hd__o221a_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ _13885_/Q _08363_/X _08126_/X _08364_/X _08359_/X vssd1 vssd1 vccd1 vccd1
+ _13885_/D sky130_fd_sc_hd__o221a_1
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07317_ _07714_/A vssd1 vssd1 vccd1 vccd1 _07317_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08297_ _08329_/A vssd1 vssd1 vccd1 vccd1 _08297_/X sky130_fd_sc_hd__buf_2
XFILLER_165_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ _07282_/A vssd1 vssd1 vccd1 vccd1 _07248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07179_ _09336_/A vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10190_ _11655_/A vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__buf_2
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12536_/X input351/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12900_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _13996_/CLK _13880_/D vssd1 vssd1 vccd1 vccd1 _13880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12831_ _12518_/X _12830_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12831_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12762_ _09556_/X _12761_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12762_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ _14621_/CLK _14501_/D vssd1 vssd1 vccd1 vccd1 _14501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _14123_/Q vssd1 vssd1 vccd1 vccd1 _11713_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12693_ _09595_/X _12692_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14527_/CLK _14432_/D vssd1 vssd1 vccd1 vccd1 _14432_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _14239_/Q _10696_/A _14434_/Q _10697_/A _11643_/X vssd1 vssd1 vccd1 vccd1
+ _11699_/B sky130_fd_sc_hd__a221oi_2
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14363_ _14633_/CLK _14363_/D vssd1 vssd1 vccd1 vccd1 _14363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 io_in[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
X_11575_ _11573_/Y _11439_/X _11574_/Y _11441_/X vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 io_in[33] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XFILLER_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 io_in[9] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_1
XFILLER_196_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13314_ _14538_/CLK _13314_/D vssd1 vssd1 vccd1 vccd1 _13314_/Q sky130_fd_sc_hd__dfxtp_1
X_10526_ _13389_/Q _10305_/X _13701_/Q _10440_/X vssd1 vssd1 vccd1 vccd1 _10526_/X
+ sky130_fd_sc_hd__a22o_1
Xinput49 la_data_in[109] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_183_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14294_ _14529_/CLK _14294_/D vssd1 vssd1 vccd1 vccd1 _14294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13245_ _14538_/CLK _13245_/D vssd1 vssd1 vccd1 vccd1 _13277_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10457_ _11655_/A vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _12667_/X input346/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10388_ _13387_/Q _10305_/X _13699_/Q _10173_/X vssd1 vssd1 vccd1 vccd1 _10388_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12127_ vssd1 vssd1 vccd1 vccd1 _12127_/HI _12127_/LO sky130_fd_sc_hd__conb_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater617 _13018_/S vssd1 vssd1 vccd1 vccd1 _13050_/S sky130_fd_sc_hd__buf_8
X_12058_ _12065_/A vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__buf_2
XFILLER_6_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater628 _12322_/S vssd1 vssd1 vccd1 vccd1 _12318_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_117_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater639 _14595_/CLK vssd1 vssd1 vccd1 vccd1 _14573_/CLK sky130_fd_sc_hd__buf_8
XFILLER_152_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11009_ _13991_/Q vssd1 vssd1 vccd1 vccd1 _11009_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06550_ _06853_/A _06740_/A vssd1 vssd1 vccd1 vccd1 _06743_/A sky130_fd_sc_hd__or2_2
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08220_ _13965_/Q _08211_/X _08119_/X _08213_/X _08214_/X vssd1 vssd1 vccd1 vccd1
+ _13965_/D sky130_fd_sc_hd__o221a_1
XFILLER_18_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08151_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08151_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07102_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07102_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08082_ _14020_/Q _08078_/X _07788_/X _08079_/X _08075_/X vssd1 vssd1 vccd1 vccd1
+ _14020_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07033_ _14551_/Q _07025_/X _06745_/X _07027_/X _07028_/X vssd1 vssd1 vccd1 vccd1
+ _14551_/D sky130_fd_sc_hd__o221a_1
XFILLER_200_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ _13580_/Q _08894_/A _08983_/X _08897_/A _08975_/X vssd1 vssd1 vccd1 vccd1
+ _13580_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _07935_/A vssd1 vssd1 vccd1 vccd1 _07935_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07866_ _14139_/Q _07863_/X _07784_/X _07864_/X _07865_/X vssd1 vssd1 vccd1 vccd1
+ _14139_/D sky130_fd_sc_hd__o221a_1
XFILLER_99_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09605_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__buf_4
XFILLER_95_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06817_ _08169_/A vssd1 vssd1 vccd1 vccd1 _06817_/X sky130_fd_sc_hd__buf_2
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07797_ _14173_/Q _07704_/A _07796_/X _07706_/A _07794_/X vssd1 vssd1 vccd1 vccd1
+ _14173_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09536_ _09588_/A vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__buf_2
X_06748_ _08119_/A vssd1 vssd1 vccd1 vccd1 _06748_/X sky130_fd_sc_hd__buf_2
XFILLER_38_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _13286_/Q _09464_/X _12281_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _13286_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06679_ _08979_/A _06575_/Y _06617_/Y _08983_/A vssd1 vssd1 vccd1 vccd1 _06679_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08418_ _13857_/Q _08415_/X _08199_/X _08417_/X _08406_/X vssd1 vssd1 vccd1 vccd1
+ _13857_/D sky130_fd_sc_hd__o221a_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09398_ _09401_/A _13143_/X vssd1 vssd1 vccd1 vccd1 _13336_/D sky130_fd_sc_hd__and2_1
XFILLER_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08349_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08349_/X sky130_fd_sc_hd__buf_2
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11360_ _11355_/Y _11161_/X _11356_/Y _11163_/X _11359_/X vssd1 vssd1 vccd1 vccd1
+ _11395_/A sky130_fd_sc_hd__o221a_2
XFILLER_165_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10309_/Y _10181_/X _10310_/Y _10184_/X vssd1 vssd1 vccd1 vccd1 _10311_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11291_ _11281_/Y _11176_/X _11284_/X _11287_/X _11290_/X vssd1 vssd1 vccd1 vccd1
+ _11313_/C sky130_fd_sc_hd__o2111a_4
X_13030_ _13029_/X _12594_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13030_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10242_ _10242_/A vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _10173_/A vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ _14169_/CLK _13932_/D vssd1 vssd1 vccd1 vccd1 _13932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ _14100_/CLK _13863_/D vssd1 vssd1 vccd1 vccd1 _13863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12814_ _12515_/X _12813_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux2_1
X_13794_ _14114_/CLK _13794_/D vssd1 vssd1 vccd1 vccd1 _13794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12745_ _09547_/X _12744_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _09586_/X input357/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12676_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14415_ _14470_/CLK _14415_/D vssd1 vssd1 vccd1 vccd1 _14415_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _14472_/Q vssd1 vssd1 vccd1 vccd1 _11627_/Y sky130_fd_sc_hd__inv_2
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _14495_/CLK _14346_/D vssd1 vssd1 vccd1 vccd1 _14346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11558_ _13964_/Q vssd1 vssd1 vccd1 vccd1 _11558_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _11457_/A vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14277_ _14527_/CLK _14277_/D vssd1 vssd1 vccd1 vccd1 _14277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11489_ _14352_/Q vssd1 vssd1 vccd1 vccd1 _11489_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13228_ _13352_/CLK _13228_/D vssd1 vssd1 vccd1 vccd1 _13260_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13159_ _12657_/X _13158_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13159_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07720_ _07785_/A vssd1 vssd1 vccd1 vccd1 _07772_/A sky130_fd_sc_hd__buf_4
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07651_ _14239_/Q _07644_/X _07330_/X _07646_/X _07650_/X vssd1 vssd1 vccd1 vccd1
+ _14239_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06602_ _06602_/A vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _14276_/Q _07580_/X _07336_/X _07581_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _14276_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09321_ _13395_/Q _09318_/X _08165_/A _09319_/X _09314_/X vssd1 vssd1 vccd1 vccd1
+ _13395_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06533_ _06535_/A vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__buf_4
XFILLER_90_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09252_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08203_ _08383_/A vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__buf_4
XFILLER_33_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09183_ _13474_/Q _09179_/X _08957_/X _09180_/X _09182_/X vssd1 vssd1 vccd1 vccd1
+ _13474_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08134_ _08184_/A vssd1 vssd1 vccd1 vccd1 _08134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08065_ _14030_/Q _08061_/X _07764_/X _08062_/X _08058_/X vssd1 vssd1 vccd1 vccd1
+ _14030_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07016_ _07070_/A vssd1 vssd1 vccd1 vccd1 _07017_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput206 la_oenb[1] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__buf_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput217 la_oenb[2] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_1
XPHY_7238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08967_ _08967_/A vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__buf_4
Xinput228 la_oenb[3] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_1
XPHY_7249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput239 la_oenb[4] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_1
XPHY_6515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07918_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07918_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08898_ _13616_/Q _08894_/X _08895_/X _08897_/X _08886_/X vssd1 vssd1 vccd1 vccd1
+ _13616_/D sky130_fd_sc_hd__o221a_1
XPHY_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ _14149_/Q _07845_/X _07759_/X _07846_/X _07848_/X vssd1 vssd1 vccd1 vccd1
+ _14149_/D sky130_fd_sc_hd__o221a_1
XPHY_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _13204_/Q _10775_/X _14027_/Q _10719_/X _10859_/X vssd1 vssd1 vccd1 vccd1
+ _10860_/X sky130_fd_sc_hd__a221o_2
XFILLER_25_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _09519_/A _12400_/X vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__and2_2
XFILLER_164_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _14142_/Q vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _13370_/Q _10033_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12530_/X sky130_fd_sc_hd__mux2_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12461_ _12509_/X _06933_/Y _12461_/S vssd1 vssd1 vccd1 vccd1 _12461_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14200_ _14481_/CLK _14200_/D vssd1 vssd1 vccd1 vccd1 _14200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11412_ _11412_/A vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__buf_2
XFILLER_107_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12392_ _13207_/Q _06657_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14131_ _14173_/CLK _14131_/D vssd1 vssd1 vccd1 vccd1 _14131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11343_ _14193_/Q vssd1 vssd1 vccd1 vccd1 _11343_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14062_ _14119_/CLK _14062_/D vssd1 vssd1 vccd1 vccd1 _14062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ _13678_/Q vssd1 vssd1 vccd1 vccd1 _11274_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13013_ _12586_/X _13012_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10225_ _10212_/Y _10214_/X _10215_/Y _10217_/X _10224_/X vssd1 vssd1 vccd1 vccd1
+ _10254_/B sky130_fd_sc_hd__o221a_2
XFILLER_49_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _10156_/A vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10087_ _10099_/A _10130_/A vssd1 vssd1 vccd1 vccd1 _12485_/S sky130_fd_sc_hd__or2_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ _14146_/CLK _13915_/D vssd1 vssd1 vccd1 vccd1 _13915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13846_ _14094_/CLK _13846_/D vssd1 vssd1 vccd1 vccd1 _13846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13777_ _14130_/CLK _13777_/D vssd1 vssd1 vccd1 vccd1 _13777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10989_ _11461_/A vssd1 vssd1 vccd1 vccd1 _10989_/X sky130_fd_sc_hd__buf_1
XFILLER_204_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12728_ _09578_/X input360/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12728_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _13347_/Q _12658_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12659_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14329_ _14637_/CLK _14329_/D vssd1 vssd1 vccd1 vccd1 _14329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _13298_/Q vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__inv_2
XFILLER_28_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08821_ _13655_/Q _08818_/X _08589_/X _08820_/X _08808_/X vssd1 vssd1 vccd1 vccd1
+ _13655_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08752_ _13694_/Q _08748_/X _08589_/X _08750_/X _08751_/X vssd1 vssd1 vccd1 vccd1
+ _13694_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07703_ _07783_/A vssd1 vssd1 vccd1 vccd1 _07704_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08683_ _13730_/Q _08677_/X _08494_/X _08679_/X _08671_/X vssd1 vssd1 vccd1 vccd1
+ _13730_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _07634_/A vssd1 vssd1 vccd1 vccd1 _07634_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07565_ _14285_/Q _07561_/X _07311_/X _07563_/X _07550_/X vssd1 vssd1 vccd1 vccd1
+ _14285_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _13406_/Q _09302_/X _08137_/A _09303_/X _09298_/X vssd1 vssd1 vccd1 vccd1
+ _13406_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06516_ _12396_/S vssd1 vssd1 vccd1 vccd1 _06853_/A sky130_fd_sc_hd__inv_2
X_07496_ _14322_/Q _07488_/X _07315_/X _07490_/X _07493_/X vssd1 vssd1 vccd1 vccd1
+ _14322_/D sky130_fd_sc_hd__o221a_1
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09235_ _13445_/Q _09233_/X _08930_/X _09234_/X _09228_/X vssd1 vssd1 vccd1 vccd1
+ _13445_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09166_ _13484_/Q _09163_/X _08930_/X _09164_/X _09165_/X vssd1 vssd1 vccd1 vccd1
+ _13484_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08117_ _08117_/A vssd1 vssd1 vccd1 vccd1 _08117_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09097_ _13523_/Q _09095_/X _08930_/X _09096_/X _09093_/X vssd1 vssd1 vccd1 vccd1
+ _13523_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08048_ _14041_/Q _08045_/X _07736_/X _08046_/X _08042_/X vssd1 vssd1 vccd1 vccd1
+ _14041_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10010_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10011_/B sky130_fd_sc_hd__inv_2
XPHY_7013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__inv_2
XFILLER_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _13856_/Q vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__inv_2
XPHY_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _14178_/CLK _13700_/D vssd1 vssd1 vccd1 vccd1 _13700_/Q sky130_fd_sc_hd__dfxtp_1
X_10912_ _10910_/Y _10739_/X _10911_/Y _10741_/X vssd1 vssd1 vccd1 vccd1 _10912_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11892_ _11890_/Y _10220_/A _11891_/Y _10223_/A vssd1 vssd1 vccd1 vccd1 _11892_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13631_ _14071_/CLK _13631_/D vssd1 vssd1 vccd1 vccd1 _13631_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _13630_/Q vssd1 vssd1 vccd1 vccd1 _10843_/Y sky130_fd_sc_hd__inv_2
XPHY_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13562_ _14114_/CLK _13562_/D vssd1 vssd1 vccd1 vccd1 _13562_/Q sky130_fd_sc_hd__dfxtp_1
X_10774_ _10764_/Y _10702_/X _10767_/X _10770_/X _10773_/X vssd1 vssd1 vccd1 vccd1
+ _10797_/C sky130_fd_sc_hd__o2111a_4
XFILLER_164_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _13356_/Q _10054_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12513_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13493_ _14481_/CLK _13493_/D vssd1 vssd1 vccd1 vccd1 _13493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12444_ _12443_/X _06912_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12375_ _13213_/Q _12374_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14114_ _14114_/CLK _14114_/D vssd1 vssd1 vccd1 vccd1 _14114_/Q sky130_fd_sc_hd__dfxtp_1
X_11326_ _13842_/Q vssd1 vssd1 vccd1 vccd1 _11326_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14045_ _14047_/CLK _14045_/D vssd1 vssd1 vccd1 vccd1 _14045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11257_ _11252_/Y _11199_/X _11253_/Y _11201_/X _11256_/X vssd1 vssd1 vccd1 vccd1
+ _11270_/B sky130_fd_sc_hd__o221a_1
XFILLER_84_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _11665_/A vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11188_ _11424_/A vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ _10146_/A _12430_/X vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ _14107_/CLK _13829_/D vssd1 vssd1 vccd1 vccd1 _13829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07350_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07350_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_206_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07281_ _14418_/Q _07274_/X _06801_/X _07275_/X _07279_/X vssd1 vssd1 vccd1 vccd1
+ _14418_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09020_ _13564_/Q _09014_/X _08925_/X _09015_/X _09019_/X vssd1 vssd1 vccd1 vccd1
+ _13564_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09922_ _13316_/Q vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__inv_2
XFILLER_119_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _09853_/A vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08804_ _13663_/Q _08800_/X _08648_/X _08801_/X _08802_/X vssd1 vssd1 vccd1 vccd1
+ _13663_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09784_ _09784_/A _09843_/A vssd1 vssd1 vccd1 vccd1 _09785_/B sky130_fd_sc_hd__or2_2
XFILLER_45_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06996_ _14562_/Q vssd1 vssd1 vccd1 vccd1 _06996_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08735_ _13700_/Q _08730_/X _08572_/X _08731_/X _08728_/X vssd1 vssd1 vccd1 vccd1
+ _13700_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_108 _10475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08666_ _13739_/Q _08662_/X _08490_/X _08663_/X _08665_/X vssd1 vssd1 vccd1 vccd1
+ _13739_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 _10838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07617_/A vssd1 vssd1 vccd1 vccd1 _07617_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08597_ _13775_/Q _08588_/X _08496_/X _08591_/X _08592_/X vssd1 vssd1 vccd1 vccd1
+ _13775_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _14291_/Q _07541_/X _07396_/X _07542_/X _07544_/X vssd1 vssd1 vccd1 vccd1
+ _14291_/D sky130_fd_sc_hd__o221a_1
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07479_ _14327_/Q _07411_/A _07403_/X _07414_/A _07476_/X vssd1 vssd1 vccd1 vccd1
+ _14327_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _13455_/Q _09215_/X _07719_/A _09217_/X _09209_/X vssd1 vssd1 vccd1 vccd1
+ _13455_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ _14292_/Q vssd1 vssd1 vccd1 vccd1 _10490_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ _09173_/A vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12160_ vssd1 vssd1 vccd1 vccd1 _12160_/HI _12160_/LO sky130_fd_sc_hd__conb_1
XFILLER_159_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ _13915_/Q vssd1 vssd1 vccd1 vccd1 _11111_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12091_ vssd1 vssd1 vccd1 vccd1 _12091_/HI _12091_/LO sky130_fd_sc_hd__conb_1
XFILLER_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ _11042_/A vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12576_/X _12992_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _14479_/Q vssd1 vssd1 vccd1 vccd1 _11944_/Y sky130_fd_sc_hd__inv_2
XPHY_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11875_ _13971_/Q vssd1 vssd1 vccd1 vccd1 _11875_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ _14173_/CLK _13614_/D vssd1 vssd1 vccd1 vccd1 _13614_/Q sky130_fd_sc_hd__dfxtp_1
X_10826_ _14299_/Q vssd1 vssd1 vccd1 vccd1 _10826_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14594_ _14595_/CLK _14594_/D vssd1 vssd1 vccd1 vccd1 _14594_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13545_ _14121_/CLK _13545_/D vssd1 vssd1 vccd1 vccd1 _13545_/Q sky130_fd_sc_hd__dfxtp_1
X_10757_ _13433_/Q vssd1 vssd1 vccd1 vccd1 _10757_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13476_ _14188_/CLK _13476_/D vssd1 vssd1 vccd1 vccd1 _13476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10688_ _13432_/Q vssd1 vssd1 vccd1 vccd1 _10688_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12427_ _12426_/X _06886_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12427_/X sky130_fd_sc_hd__mux2_1
X_12358_ _12357_/X _13203_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12358_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11309_ _14465_/Q vssd1 vssd1 vccd1 vccd1 _11309_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12289_ _11823_/Y _14554_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12289_/X sky130_fd_sc_hd__mux2_4
XFILLER_99_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14028_ _14119_/CLK _14028_/D vssd1 vssd1 vccd1 vccd1 _14028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06850_ _12396_/S _06850_/B vssd1 vssd1 vccd1 vccd1 _06850_/X sky130_fd_sc_hd__and2_1
XFILLER_56_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06781_ _08144_/A vssd1 vssd1 vccd1 vccd1 _06781_/X sky130_fd_sc_hd__buf_2
XFILLER_83_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _13806_/Q _08513_/X _08519_/X _08515_/X _08511_/X vssd1 vssd1 vccd1 vccd1
+ _13806_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08451_ _13838_/Q _08444_/X _08146_/X _08445_/X _08449_/X vssd1 vssd1 vccd1 vccd1
+ _13838_/D sky130_fd_sc_hd__o221a_1
XFILLER_184_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07402_ _14367_/Q _07307_/A _07401_/X _07309_/A _07397_/X vssd1 vssd1 vccd1 vccd1
+ _14367_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _13875_/Q _08379_/X _08153_/X _08380_/X _08375_/X vssd1 vssd1 vccd1 vccd1
+ _13875_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07333_ _07371_/A vssd1 vssd1 vccd1 vccd1 _07333_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07264_ _14428_/Q _07257_/X _06766_/X _07258_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _14428_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09003_ _09048_/A vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__buf_2
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07195_ _14466_/Q _07193_/X _06771_/X _07194_/X _07189_/X vssd1 vssd1 vccd1 vccd1
+ _14466_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09905_ _09905_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__or2_1
XFILLER_173_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09836_ _13328_/Q _09833_/Y _09779_/B vssd1 vssd1 vccd1 vccd1 _09836_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06979_ _14567_/Q vssd1 vssd1 vccd1 vccd1 _06979_/Y sky130_fd_sc_hd__inv_2
X_09767_ _13321_/Q vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__inv_2
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _13711_/Q _08714_/X _08546_/X _08715_/X _08712_/X vssd1 vssd1 vccd1 vccd1
+ _13711_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _09726_/A vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08649_ _13748_/Q _08643_/X _08648_/X _08644_/X _08646_/X vssd1 vssd1 vccd1 vccd1
+ _13748_/D sky130_fd_sc_hd__o221a_1
XPHY_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11660_/A vssd1 vssd1 vccd1 vccd1 _11660_/X sky130_fd_sc_hd__clkbuf_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10611_ _14217_/Q _10437_/X _14412_/Q _10438_/X _10610_/X vssd1 vssd1 vccd1 vccd1
+ _10644_/B sky130_fd_sc_hd__a221oi_2
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11591_ _14082_/Q vssd1 vssd1 vccd1 vccd1 _11591_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13330_ _14639_/CLK _13330_/D vssd1 vssd1 vccd1 vccd1 _13330_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10542_ _14488_/Q vssd1 vssd1 vccd1 vccd1 _10542_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13261_ _14639_/CLK _13261_/D vssd1 vssd1 vccd1 vccd1 _13261_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10473_ _11431_/A vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__clkbuf_1
X_13192_ _14071_/CLK _13192_/D vssd1 vssd1 vccd1 vccd1 _13192_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12143_ vssd1 vssd1 vccd1 vccd1 _12143_/HI _12143_/LO sky130_fd_sc_hd__conb_1
XFILLER_139_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12074_ _06492_/Y _09460_/X _09513_/B _07004_/A vssd1 vssd1 vccd1 vccd1 _14639_/D
+ sky130_fd_sc_hd__a31oi_2
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11025_ _14264_/Q vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12568_/X input331/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__mux2_1
XPHY_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11927_ _13575_/Q _10206_/A _13816_/Q _10209_/A vssd1 vssd1 vccd1 vccd1 _11927_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11858_ _11853_/Y _11679_/X _11854_/Y _11681_/X _11857_/X vssd1 vssd1 vccd1 vccd1
+ _11865_/C sky130_fd_sc_hd__o221a_1
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_19 _11907_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10809_ _13870_/Q vssd1 vssd1 vccd1 vccd1 _10809_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ _14242_/Q _11406_/A _14437_/Q _11407_/A vssd1 vssd1 vccd1 vccd1 _11789_/X
+ sky130_fd_sc_hd__a22o_2
X_14577_ _14595_/CLK _14577_/D vssd1 vssd1 vccd1 vccd1 _14577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _14120_/CLK _13528_/D vssd1 vssd1 vccd1 vccd1 _13528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13459_ _14169_/CLK _13459_/D vssd1 vssd1 vccd1 vccd1 _13459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _08411_/A _08890_/B _08584_/C _08091_/D vssd1 vssd1 vccd1 vccd1 _11633_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06902_ _14588_/Q vssd1 vssd1 vccd1 vccd1 _06902_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07882_ _07882_/A vssd1 vssd1 vccd1 vccd1 _07882_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06833_ _08977_/A vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09621_ _14596_/Q _14592_/Q _06869_/X _06886_/Y vssd1 vssd1 vccd1 vccd1 _09621_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09560_/A _12388_/X vssd1 vssd1 vccd1 vccd1 _09552_/X sky130_fd_sc_hd__and2_1
XFILLER_42_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06764_ _14624_/Q _06751_/X _06763_/X _06754_/X _06749_/X vssd1 vssd1 vccd1 vccd1
+ _14624_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08503_ _08554_/A vssd1 vssd1 vccd1 vccd1 _08503_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _13274_/Q _09479_/X _12269_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _13274_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06695_ _06662_/X _06694_/Y _06662_/X _06694_/Y vssd1 vssd1 vccd1 vccd1 _06695_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08434_ _13849_/Q _08425_/X _08117_/X _08427_/X _08433_/X vssd1 vssd1 vccd1 vccd1
+ _13849_/D sky130_fd_sc_hd__o221a_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ _13886_/Q _08363_/X _08123_/X _08364_/X _08359_/X vssd1 vssd1 vccd1 vccd1
+ _13886_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07316_ _14400_/Q _07307_/X _07315_/X _07309_/X _07301_/X vssd1 vssd1 vccd1 vccd1
+ _14400_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08296_ _08383_/A vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ _07290_/A vssd1 vssd1 vccd1 vccd1 _07282_/A sky130_fd_sc_hd__buf_4
XFILLER_30_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07178_ _14475_/Q _07174_/X _06738_/X _07176_/X _07169_/X vssd1 vssd1 vccd1 vccd1
+ _14475_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _13350_/Q _09816_/Y _09818_/Y _09816_/A vssd1 vssd1 vccd1 vccd1 _09819_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12830_ _12518_/X _12829_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12761_ _09556_/X _12760_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14500_ _14621_/CLK _14500_/D vssd1 vssd1 vccd1 vccd1 _14500_/Q sky130_fd_sc_hd__dfxtp_1
X_11712_ _13850_/Q vssd1 vssd1 vccd1 vccd1 _11712_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12692_ _09595_/X input341/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11643_ _13413_/Q _11514_/X _13725_/Q _11642_/X vssd1 vssd1 vccd1 vccd1 _11643_/X
+ sky130_fd_sc_hd__a22o_2
X_14431_ _14611_/CLK _14431_/D vssd1 vssd1 vccd1 vccd1 _14431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _14633_/CLK _14362_/D vssd1 vssd1 vccd1 vccd1 _14362_/Q sky130_fd_sc_hd__dfxtp_1
X_11574_ _14393_/Q vssd1 vssd1 vccd1 vccd1 _11574_/Y sky130_fd_sc_hd__inv_2
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 io_in[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XFILLER_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 io_in[34] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10525_ _10520_/Y _10425_/X _10521_/Y _10428_/X _10524_/X vssd1 vssd1 vccd1 vccd1
+ _10561_/A sky130_fd_sc_hd__o221a_2
Xinput39 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_6
X_13313_ _14573_/CLK _13313_/D vssd1 vssd1 vccd1 vccd1 _13313_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14293_ _14529_/CLK _14293_/D vssd1 vssd1 vccd1 vccd1 _14293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13244_ _13368_/CLK _13244_/D vssd1 vssd1 vccd1 vccd1 _13276_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10456_ _14097_/Q vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13175_ _12665_/X _13174_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__mux2_1
X_10387_ _10382_/Y _10150_/X _10383_/Y _10153_/X _10386_/X vssd1 vssd1 vccd1 vccd1
+ _10422_/A sky130_fd_sc_hd__o221a_2
XFILLER_151_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12126_ vssd1 vssd1 vccd1 vccd1 _12126_/HI _12126_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12057_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__buf_2
XFILLER_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater618 _13018_/S vssd1 vssd1 vccd1 vccd1 _12954_/S sky130_fd_sc_hd__buf_8
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater629 _10111_/A vssd1 vssd1 vccd1 vccd1 _10114_/A sky130_fd_sc_hd__buf_8
XFILLER_93_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11008_ _11006_/Y _10947_/X _11007_/Y _10949_/X vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12558_/X _12958_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12959_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14629_ _14629_/CLK _14629_/D vssd1 vssd1 vccd1 vccd1 _14629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08150_ _08150_/A vssd1 vssd1 vccd1 vccd1 _08150_/X sky130_fd_sc_hd__buf_4
XFILLER_144_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07101_ _07144_/A vssd1 vssd1 vccd1 vccd1 _07136_/A sky130_fd_sc_hd__buf_4
XFILLER_105_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08081_ _14021_/Q _08078_/X _07867_/X _08079_/X _08075_/X vssd1 vssd1 vccd1 vccd1
+ _14021_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ _14552_/Q _07025_/X _07031_/X _07027_/X _07028_/X vssd1 vssd1 vccd1 vccd1
+ _14552_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08983_ _08983_/A vssd1 vssd1 vccd1 vccd1 _08983_/X sky130_fd_sc_hd__buf_4
XFILLER_142_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07934_ _07934_/A vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07865_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07865_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09604_/A vssd1 vssd1 vccd1 vccd1 _12064_/A sky130_fd_sc_hd__buf_4
X_06816_ _08965_/A vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07796_ _08186_/A vssd1 vssd1 vccd1 vccd1 _07796_/X sky130_fd_sc_hd__buf_4
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06747_ _08914_/A vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09535_ _09535_/A vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__buf_2
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09480_/A vssd1 vssd1 vccd1 vccd1 _09466_/X sky130_fd_sc_hd__clkbuf_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06678_ _06675_/X _06677_/X _06675_/X _06677_/X vssd1 vssd1 vccd1 vccd1 _06678_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08417_ _08417_/A vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ _09401_/A _13139_/X vssd1 vssd1 vccd1 vccd1 _13337_/D sky130_fd_sc_hd__and2_1
XFILLER_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08348_ _13895_/Q _08344_/X _08099_/X _08346_/X _08336_/X vssd1 vssd1 vccd1 vccd1
+ _13895_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08279_ _13934_/Q _08274_/X _08099_/X _08276_/X _08278_/X vssd1 vssd1 vccd1 vccd1
+ _13934_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10310_ _13860_/Q vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11290_ _11288_/Y _11188_/X _11289_/Y _11190_/X vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10241_ _11689_/A vssd1 vssd1 vccd1 vccd1 _10242_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ _11642_/A vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__buf_4
XFILLER_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput490 _12122_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13931_ _14169_/CLK _13931_/D vssd1 vssd1 vccd1 vccd1 _13931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13862_ _14100_/CLK _13862_/D vssd1 vssd1 vccd1 vccd1 _13862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12813_ _12515_/X _12812_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12813_/X sky130_fd_sc_hd__mux2_1
X_13793_ _14120_/CLK _13793_/D vssd1 vssd1 vccd1 vccd1 _13793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12744_ _09547_/X input342/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12744_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12675_ _09582_/X _12674_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13197_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14414_ _14470_/CLK _14414_/D vssd1 vssd1 vccd1 vccd1 _14414_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _13490_/Q vssd1 vssd1 vccd1 vccd1 _11626_/Y sky130_fd_sc_hd__inv_2
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ _14627_/CLK _14345_/D vssd1 vssd1 vccd1 vccd1 _14345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11557_ _14237_/Q _11406_/X _14432_/Q _11407_/X _11556_/X vssd1 vssd1 vccd1 vccd1
+ _11590_/B sky130_fd_sc_hd__a221oi_2
XFILLER_89_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _11691_/A vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__buf_4
XFILLER_32_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14276_ _14527_/CLK _14276_/D vssd1 vssd1 vccd1 vccd1 _14276_/Q sky130_fd_sc_hd__dfxtp_1
X_11488_ _14508_/Q vssd1 vssd1 vccd1 vccd1 _11488_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10439_ _11642_/A vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13227_ _13352_/CLK _13227_/D vssd1 vssd1 vccd1 vccd1 _13259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_119_1914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13158_ _13157_/X _12657_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12109_ vssd1 vssd1 vccd1 vccd1 _12109_/HI _12109_/LO sky130_fd_sc_hd__conb_1
X_13089_ _12623_/X _13088_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07650_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07650_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06601_ _06603_/A vssd1 vssd1 vccd1 vccd1 _08957_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _07606_/A vssd1 vssd1 vccd1 vccd1 _07581_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09320_ _13396_/Q _09318_/X _08162_/A _09319_/X _09314_/X vssd1 vssd1 vccd1 vccd1
+ _13396_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06532_ _06532_/A vssd1 vssd1 vccd1 vccd1 _06532_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _13435_/Q _09249_/X _08957_/X _09250_/X _09244_/X vssd1 vssd1 vccd1 vccd1
+ _13435_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08202_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_178_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09182_ _09219_/A vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08133_ _08133_/A vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__buf_4
XFILLER_175_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08064_ _14031_/Q _08061_/X _07762_/X _08062_/X _08058_/X vssd1 vssd1 vccd1 vccd1
+ _14031_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07015_ _07809_/A vssd1 vssd1 vccd1 vccd1 _07015_/X sky130_fd_sc_hd__buf_2
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput207 la_oenb[20] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_1
XPHY_7228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput218 la_oenb[30] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_1
XPHY_7239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08966_ _13588_/Q _08956_/X _08965_/X _08958_/X _08963_/X vssd1 vssd1 vccd1 vccd1
+ _13588_/D sky130_fd_sc_hd__o221a_1
Xinput229 la_oenb[40] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_1
XPHY_6505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07917_ _14111_/Q _07910_/X _07755_/X _07911_/X _07913_/X vssd1 vssd1 vccd1 vccd1
+ _14111_/D sky130_fd_sc_hd__o221a_1
XPHY_6538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08897_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08897_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _07886_/A vssd1 vssd1 vccd1 vccd1 _07848_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07779_ _14180_/Q _07770_/X _07778_/X _07772_/X _07768_/X vssd1 vssd1 vccd1 vccd1
+ _14180_/D sky130_fd_sc_hd__o221a_1
X_09518_ _09509_/X _09514_/X _13286_/Q _09517_/X vssd1 vssd1 vccd1 vccd1 _13254_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _13908_/Q vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09450_/A _12927_/X vssd1 vssd1 vccd1 vccd1 _13294_/D sky130_fd_sc_hd__and2_1
XFILLER_129_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12459_/X _06930_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11411_ _13961_/Q vssd1 vssd1 vccd1 vccd1 _11411_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12391_ _12390_/X _13208_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _14130_/CLK _14130_/D vssd1 vssd1 vccd1 vccd1 _14130_/Q sky130_fd_sc_hd__dfxtp_1
X_11342_ _13601_/Q vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ _14139_/CLK _14061_/D vssd1 vssd1 vccd1 vccd1 _14061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ _13444_/Q vssd1 vssd1 vccd1 vccd1 _11273_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10224_ _10218_/Y _10220_/X _10221_/Y _10223_/X vssd1 vssd1 vccd1 vccd1 _10224_/X
+ sky130_fd_sc_hd__o22a_1
X_13012_ _12586_/X input338/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10155_ _11637_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10086_ _10098_/A _10122_/A vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__or2_1
XFILLER_188_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13914_ _14146_/CLK _13914_/D vssd1 vssd1 vccd1 vccd1 _13914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13845_ _14110_/CLK _13845_/D vssd1 vssd1 vccd1 vccd1 _13845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13776_ _14130_/CLK _13776_/D vssd1 vssd1 vccd1 vccd1 _13776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _14458_/Q vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12727_ _09576_/X _12726_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13200_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _09810_/Y _13347_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _11599_/Y _11412_/X _11602_/X _11605_/X _11608_/X vssd1 vssd1 vccd1 vccd1
+ _11631_/C sky130_fd_sc_hd__o2111a_4
XFILLER_89_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12589_ _09930_/X _13318_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14328_ _14637_/CLK _14328_/D vssd1 vssd1 vccd1 vccd1 _14328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14259_ _14305_/CLK _14259_/D vssd1 vssd1 vccd1 vccd1 _14259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08820_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08751_ _08777_/A vssd1 vssd1 vccd1 vccd1 _08751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07702_ _07785_/A vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__inv_2
X_08682_ _13731_/Q _08677_/X _08492_/X _08679_/X _08671_/X vssd1 vssd1 vccd1 vccd1
+ _13731_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07633_ _07687_/A vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _14286_/Q _07561_/X _07412_/X _07563_/X _07550_/X vssd1 vssd1 vccd1 vccd1
+ _14286_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06515_ _06515_/A1 _06492_/Y _09512_/A _06514_/X vssd1 vssd1 vccd1 vccd1 _14638_/D
+ sky130_fd_sc_hd__o22ai_4
XFILLER_55_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09303_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07495_ _14323_/Q _07488_/X _07313_/X _07490_/X _07493_/X vssd1 vssd1 vccd1 vccd1
+ _14323_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09234_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09234_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ _09173_/A vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ _14006_/Q _08109_/X _07825_/X _08112_/X _08106_/X vssd1 vssd1 vccd1 vccd1
+ _14006_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09096_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08047_ _14042_/Q _08045_/X _07733_/X _08046_/X _08042_/X vssd1 vssd1 vccd1 vccd1
+ _14042_/D sky130_fd_sc_hd__o221a_1
XFILLER_102_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09998_ _13370_/Q _09998_/B vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__nand2_1
XPHY_7036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08949_ _13595_/Q _08944_/X _08948_/X _08946_/X _08938_/X vssd1 vssd1 vccd1 vccd1
+ _13595_/D sky130_fd_sc_hd__o221a_1
XPHY_6335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _11958_/Y _10181_/A _11959_/Y _10184_/A vssd1 vssd1 vccd1 vccd1 _11960_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10911_ _14262_/Q vssd1 vssd1 vccd1 vccd1 _10911_/Y sky130_fd_sc_hd__inv_2
XPHY_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11891_ _14400_/Q vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__inv_2
XPHY_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _14071_/CLK _13630_/D vssd1 vssd1 vccd1 vccd1 _13630_/Q sky130_fd_sc_hd__dfxtp_1
X_10842_ _13669_/Q vssd1 vssd1 vccd1 vccd1 _10842_/Y sky130_fd_sc_hd__inv_2
XPHY_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13561_ _14114_/CLK _13561_/D vssd1 vssd1 vccd1 vccd1 _13561_/Q sky130_fd_sc_hd__dfxtp_1
X_10773_ _10771_/Y _10714_/X _10772_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _10773_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12512_ _13357_/Q _10055_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12512_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13492_ _14481_/CLK _13492_/D vssd1 vssd1 vccd1 vccd1 _13492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12443_ _12509_/X _06912_/Y _12443_/S vssd1 vssd1 vccd1 vccd1 _12443_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12374_ _13213_/Q _06609_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14113_ _14114_/CLK _14113_/D vssd1 vssd1 vccd1 vccd1 _14113_/Q sky130_fd_sc_hd__dfxtp_1
X_11325_ _11323_/Y _11178_/X _11324_/Y _11180_/X vssd1 vssd1 vccd1 vccd1 _11325_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14044_ _14047_/CLK _14044_/D vssd1 vssd1 vccd1 vccd1 _14044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ _11254_/Y _11203_/X _11255_/Y _11205_/X vssd1 vssd1 vccd1 vccd1 _11256_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _10207_/A vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__inv_2
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11187_ _13995_/Q vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10138_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _12428_/S sky130_fd_sc_hd__or2_1
XFILLER_94_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _10080_/A _12502_/X vssd1 vssd1 vccd1 vccd1 _12235_/A sky130_fd_sc_hd__nor2_8
XFILLER_97_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13828_ _14107_/CLK _13828_/D vssd1 vssd1 vccd1 vccd1 _13828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13877_/CLK _13759_/D vssd1 vssd1 vccd1 vccd1 _13759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ _14419_/Q _07274_/X _07058_/X _07275_/X _07279_/X vssd1 vssd1 vccd1 vccd1
+ _14419_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09921_ _09919_/A _09919_/B _09920_/Y vssd1 vssd1 vccd1 vccd1 _09921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09852_ _13323_/Q _09850_/Y _09774_/B vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08803_ _13664_/Q _08800_/X _08566_/X _08801_/X _08802_/X vssd1 vssd1 vccd1 vccd1
+ _13664_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09783_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__or2_1
XFILLER_80_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06995_ _07004_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _14563_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08734_ _13701_/Q _08730_/X _08570_/X _08731_/X _08728_/X vssd1 vssd1 vccd1 vccd1
+ _13701_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08665_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08665_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_109 _11447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07616_ _14255_/Q _07613_/X _07471_/X _07614_/X _07609_/X vssd1 vssd1 vccd1 vccd1
+ _14255_/D sky130_fd_sc_hd__o221a_1
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08596_ _13776_/Q _08588_/X _08494_/X _08591_/X _08592_/X vssd1 vssd1 vccd1 vccd1
+ _13776_/D sky130_fd_sc_hd__o221a_1
XPHY_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ _14292_/Q _07541_/X _07394_/X _07542_/X _07544_/X vssd1 vssd1 vccd1 vccd1
+ _14292_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07478_ _14328_/Q _07411_/A _07401_/X _07414_/A _07476_/X vssd1 vssd1 vccd1 vccd1
+ _14328_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09217_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09217_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09148_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09079_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _11105_/Y _10973_/X _11106_/Y _10975_/X _11109_/X vssd1 vssd1 vccd1 vccd1
+ _11117_/C sky130_fd_sc_hd__o221a_1
XFILLER_85_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12090_ vssd1 vssd1 vccd1 vccd1 _12090_/HI _12090_/LO sky130_fd_sc_hd__conb_1
XFILLER_46_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11041_ _11036_/Y _10923_/X _11037_/Y _10925_/X _11040_/X vssd1 vssd1 vccd1 vccd1
+ _11077_/A sky130_fd_sc_hd__o221a_4
XFILLER_81_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12992_ _12576_/X input344/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__mux2_1
XPHY_6165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11943_ _13497_/Q vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__inv_2
XPHY_6198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _13418_/Q _11747_/X _13737_/Q _12416_/S _11873_/X vssd1 vssd1 vccd1 vccd1
+ _11907_/B sky130_fd_sc_hd__a221oi_2
XPHY_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13613_ _14173_/CLK _13613_/D vssd1 vssd1 vccd1 vccd1 _13613_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _10820_/Y _10725_/X _10821_/Y _10727_/X _10824_/X vssd1 vssd1 vccd1 vccd1
+ _10838_/B sky130_fd_sc_hd__o221a_4
XFILLER_44_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14621_/CLK _14593_/D vssd1 vssd1 vccd1 vccd1 _14593_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13544_ _14121_/CLK _13544_/D vssd1 vssd1 vccd1 vccd1 _13544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10756_ _14064_/Q vssd1 vssd1 vccd1 vccd1 _10756_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13475_ _14188_/CLK _13475_/D vssd1 vssd1 vccd1 vccd1 _13475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _11397_/A vssd1 vssd1 vccd1 vccd1 _10687_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12426_ _12425_/X _06886_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12357_ _13203_/Q _12356_/X input78/X vssd1 vssd1 vccd1 vccd1 _12357_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11308_ _13483_/Q vssd1 vssd1 vccd1 vccd1 _11308_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12288_ _11866_/Y _14555_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__mux2_4
XFILLER_9_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14027_ _14120_/CLK _14027_/D vssd1 vssd1 vccd1 vccd1 _14027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11239_ _13762_/Q vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06780_ _08940_/A vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__buf_4
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _13839_/Q _08444_/X _08144_/X _08445_/X _08449_/X vssd1 vssd1 vccd1 vccd1
+ _13839_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ _08188_/A vssd1 vssd1 vccd1 vccd1 _07401_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_205_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08381_ _13876_/Q _08379_/X _08150_/X _08380_/X _08375_/X vssd1 vssd1 vccd1 vccd1
+ _13876_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07332_ _08119_/A vssd1 vssd1 vccd1 vccd1 _07332_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07263_ _14429_/Q _07257_/X _06763_/X _07258_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _14429_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09002_ _13573_/Q _08993_/X _08829_/X _08995_/X _09000_/X vssd1 vssd1 vccd1 vccd1
+ _13573_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07194_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _09904_/A _09940_/A vssd1 vssd1 vccd1 vccd1 _09905_/B sky130_fd_sc_hd__or2_1
XFILLER_154_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ _09847_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _13112_/S sky130_fd_sc_hd__and2_4
XFILLER_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09766_ _13322_/Q vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__inv_2
X_06978_ _06991_/A _06978_/B vssd1 vssd1 vccd1 vccd1 _14568_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _13712_/Q _08714_/X _08544_/X _08715_/X _08712_/X vssd1 vssd1 vccd1 vccd1
+ _13712_/D sky130_fd_sc_hd__o221a_1
XPHY_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09732_/A _10077_/A vssd1 vssd1 vccd1 vccd1 _12510_/S sky130_fd_sc_hd__nand2_4
XPHY_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _09051_/A vssd1 vssd1 vccd1 vccd1 _08648_/X sky130_fd_sc_hd__clkbuf_4
XPHY_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _08983_/A vssd1 vssd1 vccd1 vccd1 _08579_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_109_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10610_ _13391_/Q _10568_/X _13703_/Q _10440_/X vssd1 vssd1 vccd1 vccd1 _10610_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _11590_/A _11590_/B _11590_/C _11590_/D vssd1 vssd1 vccd1 vccd1 _11590_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10541_ _13197_/Q _10539_/X _14020_/Q _10469_/X _10540_/X vssd1 vssd1 vccd1 vccd1
+ _10541_/X sky130_fd_sc_hd__a221o_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13260_ _14639_/CLK _13260_/D vssd1 vssd1 vccd1 vccd1 _13260_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10472_ _11665_/A vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13191_ _14071_/CLK _13191_/D vssd1 vssd1 vccd1 vccd1 _13191_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_100_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12142_ vssd1 vssd1 vccd1 vccd1 _12142_/HI _12142_/LO sky130_fd_sc_hd__conb_1
XFILLER_124_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12073_ _09818_/Y _12035_/A _09929_/Y _09607_/A vssd1 vssd1 vccd1 vccd1 _12073_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11024_ _14186_/Q vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12975_ _12566_/X _12974_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11926_ _11916_/Y _10178_/A _11919_/X _11922_/X _11925_/X vssd1 vssd1 vccd1 vccd1
+ _11948_/C sky130_fd_sc_hd__o2111a_4
XPHY_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11855_/Y _11683_/X _11856_/Y _11685_/X vssd1 vssd1 vccd1 vccd1 _11857_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _13753_/Q vssd1 vssd1 vccd1 vccd1 _10808_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ _14621_/CLK _14576_/D vssd1 vssd1 vccd1 vccd1 _14576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11788_ _11783_/Y _11633_/X _11784_/Y _11635_/X _11787_/X vssd1 vssd1 vccd1 vccd1
+ _11823_/A sky130_fd_sc_hd__o221a_1
XFILLER_109_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13527_ _14120_/CLK _13527_/D vssd1 vssd1 vccd1 vccd1 _13527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10739_ _11449_/A vssd1 vssd1 vccd1 vccd1 _10739_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13458_ _14169_/CLK _13458_/D vssd1 vssd1 vccd1 vccd1 _13458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12409_ _12408_/X _13218_/Q _12645_/S vssd1 vssd1 vccd1 vccd1 _12409_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _14529_/CLK _13389_/D vssd1 vssd1 vccd1 vccd1 _13389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07950_ _08989_/B vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06901_ _06956_/A vssd1 vssd1 vccd1 vccd1 _06901_/X sky130_fd_sc_hd__buf_1
X_07881_ _07934_/A vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__buf_2
XFILLER_25_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ _09608_/X _09619_/X _09608_/X _09619_/X vssd1 vssd1 vccd1 vccd1 _09620_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06832_ _14605_/Q _06823_/X _06831_/X _06532_/A _06821_/X vssd1 vssd1 vccd1 vccd1
+ _14605_/D sky130_fd_sc_hd__o221a_1
XFILLER_42_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09551_ _09544_/X _09550_/X _13274_/Q _09545_/X vssd1 vssd1 vccd1 vccd1 _13242_/D
+ sky130_fd_sc_hd__o22a_1
X_06763_ _08130_/A vssd1 vssd1 vccd1 vccd1 _06763_/X sky130_fd_sc_hd__buf_2
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08502_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08554_/A sky130_fd_sc_hd__buf_2
XFILLER_97_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09482_ _13275_/Q _09479_/X _12270_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _13275_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06694_ _06670_/X _06693_/Y _06670_/X _06693_/Y vssd1 vssd1 vccd1 vccd1 _06694_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08433_ _08465_/A vssd1 vssd1 vccd1 vccd1 _08433_/X sky130_fd_sc_hd__clkbuf_2
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08364_ _08389_/A vssd1 vssd1 vccd1 vccd1 _08364_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07315_ _07712_/A vssd1 vssd1 vccd1 vccd1 _07315_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08295_ _13925_/Q _08293_/X _08123_/X _08294_/X _08288_/X vssd1 vssd1 vccd1 vccd1
+ _13925_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07246_ _14438_/Q _07238_/X _06725_/X _07240_/X _07244_/X vssd1 vssd1 vccd1 vccd1
+ _14438_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ _14476_/Q _07174_/X _06735_/X _07176_/X _07169_/X vssd1 vssd1 vccd1 vccd1
+ _14476_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09818_ _13350_/Q vssd1 vssd1 vccd1 vccd1 _09818_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09749_ _13339_/Q vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__inv_2
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _09556_/X input337/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__mux2_1
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11709_/Y _11648_/X _11710_/Y _11650_/X vssd1 vssd1 vccd1 vccd1 _11711_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12691_ _09593_/X _12690_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13193_/D sky130_fd_sc_hd__mux2_1
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14430_ _14611_/CLK _14430_/D vssd1 vssd1 vccd1 vccd1 _14430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A vssd1 vssd1 vccd1 vccd1 _11642_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _14637_/CLK _14361_/D vssd1 vssd1 vccd1 vccd1 _14361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _14627_/Q vssd1 vssd1 vccd1 vccd1 _11573_/Y sky130_fd_sc_hd__inv_2
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_in[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13312_ _14573_/CLK _13312_/D vssd1 vssd1 vccd1 vccd1 _13312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 io_in[35] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XFILLER_196_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10524_ _10522_/Y _10431_/X _10523_/Y _10434_/X vssd1 vssd1 vccd1 vccd1 _10524_/X
+ sky130_fd_sc_hd__o22a_1
X_14292_ _14529_/CLK _14292_/D vssd1 vssd1 vccd1 vccd1 _14292_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _13368_/CLK _13243_/D vssd1 vssd1 vccd1 vccd1 _13275_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_124_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10455_ _11419_/A vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13174_ _13173_/X _12665_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13174_/X sky130_fd_sc_hd__mux2_1
X_10386_ _10384_/Y _10156_/X _10385_/Y _10159_/X vssd1 vssd1 vccd1 vccd1 _10386_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ vssd1 vssd1 vccd1 vccd1 _12125_/HI _12125_/LO sky130_fd_sc_hd__conb_1
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12056_ _09787_/A _12050_/X _09899_/A _12051_/X vssd1 vssd1 vccd1 vccd1 _12056_/Y
+ sky130_fd_sc_hd__o22ai_1
Xrepeater608 _12650_/S vssd1 vssd1 vccd1 vccd1 _12634_/S sky130_fd_sc_hd__buf_8
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater619 _12974_/S vssd1 vssd1 vccd1 vccd1 _13018_/S sky130_fd_sc_hd__buf_8
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ _14108_/Q vssd1 vssd1 vccd1 vccd1 _11007_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_0_register_file.clk_i _12283_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_register_file.clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12958_ _12957_/X _12558_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11909_ _13458_/Q vssd1 vssd1 vccd1 vccd1 _11909_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12889_ _12533_/X _12888_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__mux2_1
XPHY_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ _14629_/CLK _14628_/D vssd1 vssd1 vccd1 vccd1 _14628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14559_ _14637_/CLK _14559_/D vssd1 vssd1 vccd1 vccd1 _14559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07100_ _14516_/Q _07092_/X _06725_/X _07094_/X _07096_/X vssd1 vssd1 vccd1 vccd1
+ _14516_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08080_ _14022_/Q _08078_/X _07784_/X _08079_/X _08075_/X vssd1 vssd1 vccd1 vccd1
+ _14022_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07031_ _08217_/A vssd1 vssd1 vccd1 vccd1 _07031_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08982_ _13581_/Q _08894_/A _08981_/X _08897_/A _08975_/X vssd1 vssd1 vccd1 vccd1
+ _13581_/D sky130_fd_sc_hd__o221a_1
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _14101_/Q _07926_/X _07780_/X _07927_/X _07929_/X vssd1 vssd1 vccd1 vccd1
+ _14101_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07864_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07864_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09603_ _09603_/A vssd1 vssd1 vccd1 vccd1 _12858_/S sky130_fd_sc_hd__inv_8
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06815_ _14610_/Q _06805_/X _06814_/X _06811_/X _06803_/X vssd1 vssd1 vccd1 vccd1
+ _14610_/D sky130_fd_sc_hd__o221a_1
XFILLER_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07795_ _14174_/Q _07783_/X _07792_/X _07785_/X _07794_/X vssd1 vssd1 vccd1 vccd1
+ _14174_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09534_ _09530_/X _09533_/X _13280_/Q _09531_/X vssd1 vssd1 vccd1 vccd1 _13248_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06746_ _14629_/Q _06733_/X _06745_/X _06726_/X _06730_/X vssd1 vssd1 vccd1 vccd1
+ _14629_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09465_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__buf_6
XFILLER_77_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06677_ _06571_/X _06676_/X _06571_/X _06676_/X vssd1 vssd1 vccd1 vccd1 _06677_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08416_ _08469_/A vssd1 vssd1 vccd1 vccd1 _08417_/A sky130_fd_sc_hd__clkbuf_2
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09396_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_209_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08347_ _13896_/Q _08344_/X _08199_/X _08346_/X _08336_/X vssd1 vssd1 vccd1 vccd1
+ _13896_/D sky130_fd_sc_hd__o221a_1
XFILLER_90_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _08288_/A vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__buf_2
XFILLER_192_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07229_ _14444_/Q _07164_/A _06850_/B _07166_/A _07228_/X vssd1 vssd1 vccd1 vccd1
+ _14444_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _13897_/Q vssd1 vssd1 vccd1 vccd1 _10240_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _10171_/A vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__inv_2
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput480 _12113_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput491 _12123_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13930_ _14139_/CLK _13930_/D vssd1 vssd1 vccd1 vccd1 _13930_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13861_ _14095_/CLK _13861_/D vssd1 vssd1 vccd1 vccd1 _13861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12515_/X input355/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12812_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13792_ _14120_/CLK _13792_/D vssd1 vssd1 vccd1 vccd1 _13792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12743_ _09543_/X _12742_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13212_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _09582_/X _12673_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14470_/CLK _14413_/D vssd1 vssd1 vccd1 vccd1 _14413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _14160_/Q vssd1 vssd1 vccd1 vccd1 _11625_/Y sky130_fd_sc_hd__inv_2
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14344_ _14627_/CLK _14344_/D vssd1 vssd1 vccd1 vccd1 _14344_/Q sky130_fd_sc_hd__dfxtp_1
X_11556_ _13411_/Q _11514_/X _13723_/Q _11408_/X vssd1 vssd1 vccd1 vccd1 _11556_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_102_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _14136_/Q vssd1 vssd1 vccd1 vccd1 _10507_/Y sky130_fd_sc_hd__inv_2
X_14275_ _14527_/CLK _14275_/D vssd1 vssd1 vccd1 vccd1 _14275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11487_ _13217_/Q _11485_/X _14040_/Q _11429_/X _11486_/X vssd1 vssd1 vccd1 vccd1
+ _11487_/X sky130_fd_sc_hd__a221o_4
XFILLER_13_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13226_ _13352_/CLK _13226_/D vssd1 vssd1 vccd1 vccd1 _13258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ _10697_/A vssd1 vssd1 vccd1 vccd1 _10438_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13157_ _12657_/X _13156_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
X_10369_ _13581_/Q vssd1 vssd1 vccd1 vccd1 _10369_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12108_ vssd1 vssd1 vccd1 vccd1 _12108_/HI _12108_/LO sky130_fd_sc_hd__conb_1
XFILLER_61_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088_ _12623_/X input335/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12039_ _09774_/A _12035_/X _09886_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12039_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ _06602_/A vssd1 vssd1 vccd1 vccd1 _06600_/Y sky130_fd_sc_hd__inv_2
X_07580_ _07605_/A vssd1 vssd1 vccd1 vccd1 _07580_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06531_ _06811_/A vssd1 vssd1 vccd1 vccd1 _06532_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_206_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08201_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09219_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ _08132_/A vssd1 vssd1 vccd1 vccd1 _08132_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08063_ _14032_/Q _08061_/X _07759_/X _08062_/X _08058_/X vssd1 vssd1 vccd1 vccd1
+ _14032_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07014_ _07014_/A vssd1 vssd1 vccd1 vccd1 _07014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08965_ _08965_/A vssd1 vssd1 vccd1 vccd1 _08965_/X sky130_fd_sc_hd__buf_4
Xinput208 la_oenb[21] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_1
XPHY_7229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput219 la_oenb[31] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_1
XPHY_6506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07916_ _14112_/Q _07910_/X _07753_/X _07911_/X _07913_/X vssd1 vssd1 vccd1 vccd1
+ _14112_/D sky130_fd_sc_hd__o221a_1
XPHY_6528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ _08971_/A vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__clkbuf_2
XPHY_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07847_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__buf_4
XFILLER_211_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07778_ _08169_/A vssd1 vssd1 vccd1 vccd1 _07778_/X sky130_fd_sc_hd__buf_4
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09517_ _09545_/A vssd1 vssd1 vccd1 vccd1 _09517_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06729_ _07130_/A vssd1 vssd1 vccd1 vccd1 _06785_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09450_/A _12987_/X vssd1 vssd1 vccd1 vccd1 _13295_/D sky130_fd_sc_hd__and2_1
XFILLER_164_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09379_ _09382_/A _12827_/X vssd1 vssd1 vccd1 vccd1 _13351_/D sky130_fd_sc_hd__and2_1
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11410_ _14234_/Q _11406_/X _14429_/Q _11407_/X _11409_/X vssd1 vssd1 vccd1 vccd1
+ _11465_/B sky130_fd_sc_hd__a221oi_2
XFILLER_36_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12390_ _13208_/Q _12389_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11341_ _14310_/Q vssd1 vssd1 vccd1 vccd1 _11341_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14060_ _14139_/CLK _14060_/D vssd1 vssd1 vccd1 vccd1 _14060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11272_ _14075_/Q vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13011_ _12584_/X _13010_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13011_/X sky130_fd_sc_hd__mux2_1
X_10223_ _10223_/A vssd1 vssd1 vccd1 vccd1 _10223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _13656_/Q vssd1 vssd1 vccd1 vccd1 _10154_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10085_ _10094_/A _12490_/X vssd1 vssd1 vccd1 vccd1 _12239_/A sky130_fd_sc_hd__nor2_8
XFILLER_188_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13913_ _14146_/CLK _13913_/D vssd1 vssd1 vccd1 vccd1 _13913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13844_ _14110_/CLK _13844_/D vssd1 vssd1 vccd1 vccd1 _13844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13775_ _14130_/CLK _13775_/D vssd1 vssd1 vccd1 vccd1 _13775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10987_ _11459_/A vssd1 vssd1 vccd1 vccd1 _10987_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ _09576_/X _12725_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12726_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12657_ _13348_/Q _12656_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12657_/X sky130_fd_sc_hd__mux2_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11606_/Y _11424_/X _11607_/Y _11426_/X vssd1 vssd1 vccd1 vccd1 _11608_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12588_ _13303_/Q _12587_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12588_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14327_ _14637_/CLK _14327_/D vssd1 vssd1 vccd1 vccd1 _14327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11539_ _14275_/Q vssd1 vssd1 vccd1 vccd1 _11539_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14258_ _14305_/CLK _14258_/D vssd1 vssd1 vccd1 vccd1 _14258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _13368_/CLK _13209_/D vssd1 vssd1 vccd1 vccd1 _13209_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14189_ _14305_/CLK _14189_/D vssd1 vssd1 vccd1 vccd1 _14189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08750_ _08750_/A vssd1 vssd1 vccd1 vccd1 _08750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07701_ _07952_/A _11683_/A vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__or2_2
XFILLER_22_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08681_ _13732_/Q _08677_/X _08490_/X _08679_/X _08671_/X vssd1 vssd1 vccd1 vccd1
+ _13732_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07632_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__inv_2
XFILLER_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07563_ _07563_/A vssd1 vssd1 vccd1 vccd1 _07563_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09302_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09302_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06514_ _09511_/B _06505_/X _09603_/A _09607_/A vssd1 vssd1 vccd1 vccd1 _06514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _14324_/Q _07488_/X _07311_/X _07490_/X _07493_/X vssd1 vssd1 vccd1 vccd1
+ _14324_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09164_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08115_ _14007_/Q _08109_/X _08114_/X _08112_/X _08106_/X vssd1 vssd1 vccd1 vccd1
+ _14007_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09095_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08046_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08046_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09997_ _09997_/A vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__inv_2
XPHY_7026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _08948_/A vssd1 vssd1 vccd1 vccd1 _08948_/X sky130_fd_sc_hd__buf_4
XPHY_7059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _08879_/A vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__buf_6
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10910_ _14184_/Q vssd1 vssd1 vccd1 vccd1 _10910_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _14634_/Q vssd1 vssd1 vccd1 vccd1 _11890_/Y sky130_fd_sc_hd__inv_2
XPHY_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _13435_/Q vssd1 vssd1 vccd1 vccd1 _10841_/Y sky130_fd_sc_hd__inv_2
XPHY_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13560_ _14114_/CLK _13560_/D vssd1 vssd1 vccd1 vccd1 _13560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _13511_/Q vssd1 vssd1 vccd1 vccd1 _10772_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _13358_/Q _10056_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12511_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13491_ _14481_/CLK _13491_/D vssd1 vssd1 vccd1 vccd1 _13491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12442_ _12441_/X _06909_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12442_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12373_ _12372_/X _13214_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12373_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14112_ _14114_/CLK _14112_/D vssd1 vssd1 vccd1 vccd1 _14112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11324_ _13881_/Q vssd1 vssd1 vccd1 vccd1 _11324_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14043_ _14047_/CLK _14043_/D vssd1 vssd1 vccd1 vccd1 _14043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11255_ _14386_/Q vssd1 vssd1 vccd1 vccd1 _11255_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ _10206_/A vssd1 vssd1 vccd1 vccd1 _10206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11182_/Y _11183_/X _11184_/Y _11185_/X vssd1 vssd1 vccd1 vccd1 _11186_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10137_ _10137_/A _12433_/X vssd1 vssd1 vccd1 vccd1 _10137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10068_ _10079_/A _10115_/A vssd1 vssd1 vccd1 vccd1 _12500_/S sky130_fd_sc_hd__or2_1
XPHY_6870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13827_ _14100_/CLK _13827_/D vssd1 vssd1 vccd1 vccd1 _13827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13758_ _13877_/CLK _13758_/D vssd1 vssd1 vccd1 vccd1 _13758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _09565_/X _12708_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13689_ _14139_/CLK _13689_/D vssd1 vssd1 vccd1 vccd1 _13689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _09923_/B vssd1 vssd1 vccd1 vccd1 _09920_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09851_ _09772_/A _09772_/B _09850_/Y vssd1 vssd1 vccd1 vccd1 _09851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08802_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09782_ _09782_/A _09840_/A vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__or2_2
XFILLER_189_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06994_ _06857_/A _12319_/X _06993_/Y _06861_/A vssd1 vssd1 vccd1 vccd1 _06995_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08733_ _13702_/Q _08730_/X _08648_/X _08731_/X _08728_/X vssd1 vssd1 vccd1 vccd1
+ _13702_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08664_ _13740_/Q _08662_/X _08589_/X _08663_/X _08653_/X vssd1 vssd1 vccd1 vccd1
+ _13740_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07615_ _14256_/Q _07613_/X _07388_/X _07614_/X _07609_/X vssd1 vssd1 vccd1 vccd1
+ _14256_/D sky130_fd_sc_hd__o221a_1
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08595_ _13777_/Q _08588_/X _08492_/X _08591_/X _08592_/X vssd1 vssd1 vccd1 vccd1
+ _13777_/D sky130_fd_sc_hd__o221a_1
XPHY_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _14293_/Q _07541_/X _07392_/X _07542_/X _07544_/X vssd1 vssd1 vccd1 vccd1
+ _14293_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07477_ _14329_/Q _07411_/A _07399_/X _07414_/A _07476_/X vssd1 vssd1 vccd1 vccd1
+ _14329_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09216_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__buf_6
XFILLER_91_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09147_ _09189_/A vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__buf_6
XFILLER_104_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09078_ _09120_/A vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08029_ _14051_/Q _08025_/X _07708_/X _08027_/X _08017_/X vssd1 vssd1 vccd1 vccd1
+ _14051_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11040_ _11038_/Y _10927_/X _11039_/Y _10929_/X vssd1 vssd1 vccd1 vccd1 _11040_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12574_/X _12990_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ _14167_/Q vssd1 vssd1 vccd1 vccd1 _11942_/Y sky130_fd_sc_hd__inv_2
XPHY_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11873_ _14244_/Q _11830_/X _14439_/Q _11831_/X vssd1 vssd1 vccd1 vccd1 _11873_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13612_ _14173_/CLK _13612_/D vssd1 vssd1 vccd1 vccd1 _13612_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10824_ _10822_/Y _10729_/X _10823_/Y _10731_/X vssd1 vssd1 vccd1 vccd1 _10824_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14621_/CLK _14592_/D vssd1 vssd1 vccd1 vccd1 _14592_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13543_ _14121_/CLK _13543_/D vssd1 vssd1 vccd1 vccd1 _13543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10755_ _10755_/A _10755_/B _10755_/C _10755_/D vssd1 vssd1 vccd1 vccd1 _10755_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_185_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13474_ _14146_/CLK _13474_/D vssd1 vssd1 vccd1 vccd1 _13474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10686_ _14063_/Q vssd1 vssd1 vccd1 vccd1 _10686_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12425_ _12509_/X _06886_/Y _12425_/S vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12356_ _13203_/Q _06559_/A _12368_/S vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _14153_/Q vssd1 vssd1 vccd1 vccd1 _11307_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12287_ _11907_/Y _14556_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12287_/X sky130_fd_sc_hd__mux2_4
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026_ _14120_/CLK _14026_/D vssd1 vssd1 vccd1 vccd1 _14026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11238_ _13957_/Q vssd1 vssd1 vccd1 vccd1 _11238_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11169_ _11160_/Y _11161_/X _11162_/Y _11163_/X _11168_/X vssd1 vssd1 vccd1 vccd1
+ _11229_/A sky130_fd_sc_hd__o221a_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07400_ _14368_/Q _07307_/A _07399_/X _07309_/A _07397_/X vssd1 vssd1 vccd1 vccd1
+ _14368_/D sky130_fd_sc_hd__o221a_1
XFILLER_149_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08380_ _08389_/A vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07331_ _14395_/Q _07322_/X _07330_/X _07325_/X _07319_/X vssd1 vssd1 vccd1 vccd1
+ _14395_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _07262_/A vssd1 vssd1 vccd1 vccd1 _07262_/X sky130_fd_sc_hd__buf_2
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09001_ _13574_/Q _08993_/X _08827_/X _08995_/X _09000_/X vssd1 vssd1 vccd1 vccd1
+ _13574_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07193_ _07209_/A vssd1 vssd1 vccd1 vccd1 _07193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09903_ _09903_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__or2_1
XFILLER_8_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09834_ _09777_/A _09777_/B _09833_/Y vssd1 vssd1 vccd1 vccd1 _09834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ _13323_/Q vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__inv_2
X_06977_ _06974_/X _12314_/X _06975_/Y _06976_/X vssd1 vssd1 vccd1 vccd1 _06978_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08716_ _13713_/Q _08714_/X _08541_/X _08715_/X _08712_/X vssd1 vssd1 vccd1 vccd1
+ _13713_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09696_ _09686_/X _09695_/X _09686_/X _09695_/X vssd1 vssd1 vccd1 vccd1 _10077_/A
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ _13749_/Q _08643_/X _08566_/X _08644_/X _08646_/X vssd1 vssd1 vccd1 vccd1
+ _13749_/D sky130_fd_sc_hd__o221a_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08578_ _13783_/Q _08486_/A _08577_/X _08488_/A _08575_/X vssd1 vssd1 vccd1 vccd1
+ _13783_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ _14303_/Q _07524_/X _07367_/X _07525_/X _07527_/X vssd1 vssd1 vccd1 vccd1
+ _14303_/D sky130_fd_sc_hd__o221a_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _13545_/Q _10471_/X _13786_/Q _10473_/X vssd1 vssd1 vccd1 vccd1 _10540_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _11430_/A vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12210_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ _06881_/Y _06875_/Y _06889_/Y _06886_/Y _12506_/S _12507_/S vssd1 vssd1 vccd1
+ vccd1 _13190_/X sky130_fd_sc_hd__mux4_2
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ vssd1 vssd1 vccd1 vccd1 _12141_/HI _12141_/LO sky130_fd_sc_hd__conb_1
XFILLER_178_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12072_ _09815_/A _12035_/A _09926_/A _09607_/A vssd1 vssd1 vccd1 vccd1 _12072_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_137_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11023_ _13594_/Q vssd1 vssd1 vccd1 vccd1 _11023_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12974_ _12973_/X _12566_/X _12974_/S vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__mux2_1
XPHY_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11925_ _11923_/Y _10195_/A _11924_/Y _10198_/A vssd1 vssd1 vccd1 vccd1 _11925_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11856_ _14282_/Q vssd1 vssd1 vccd1 vccd1 _11856_/Y sky130_fd_sc_hd__inv_2
XPHY_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _13948_/Q vssd1 vssd1 vccd1 vccd1 _10807_/Y sky130_fd_sc_hd__inv_2
XPHY_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _14621_/CLK _14575_/D vssd1 vssd1 vccd1 vccd1 _14575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11787_ _11785_/Y _11637_/X _11786_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _11787_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13526_ _14120_/CLK _13526_/D vssd1 vssd1 vccd1 vccd1 _13526_/Q sky130_fd_sc_hd__dfxtp_1
X_10738_ _14180_/Q vssd1 vssd1 vccd1 vccd1 _10738_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13457_ _14169_/CLK _13457_/D vssd1 vssd1 vccd1 vccd1 _13457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10669_ _14374_/Q vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12408_ _13218_/Q _12407_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _14529_/CLK _13388_/D vssd1 vssd1 vccd1 vccd1 _13388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12339_ _13193_/Q _12338_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12339_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14009_ _14094_/CLK _14009_/D vssd1 vssd1 vccd1 vccd1 _14009_/Q sky130_fd_sc_hd__dfxtp_1
X_06900_ _06918_/A vssd1 vssd1 vccd1 vccd1 _06917_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07880_ _07935_/A vssd1 vssd1 vccd1 vccd1 _07934_/A sky130_fd_sc_hd__inv_2
XFILLER_29_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06831_ _08179_/A vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09550_ _09560_/A _12385_/X vssd1 vssd1 vccd1 vccd1 _09550_/X sky130_fd_sc_hd__and2_1
XFILLER_42_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06762_ _08925_/A vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08501_ _08833_/A vssd1 vssd1 vccd1 vccd1 _08501_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ _13276_/Q _09479_/X _12271_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _13276_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06693_ _06674_/X _06692_/X _06674_/X _06692_/X vssd1 vssd1 vccd1 vccd1 _06693_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_129_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08432_ _08645_/A vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ _08388_/A vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07314_ _14401_/Q _07307_/X _07313_/X _07309_/X _07301_/X vssd1 vssd1 vccd1 vccd1
+ _14401_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08294_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07245_ _14439_/Q _07238_/X _06722_/X _07240_/X _07244_/X vssd1 vssd1 vccd1 vccd1
+ _14439_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07176_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09817_ _09815_/A _09815_/B _09816_/Y vssd1 vssd1 vccd1 vccd1 _09817_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ _13340_/Q vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__inv_2
XFILLER_21_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09679_ _09669_/X _09678_/X _09669_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _10065_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _13889_/Q vssd1 vssd1 vccd1 vccd1 _11710_/Y sky130_fd_sc_hd__inv_2
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12690_ _09593_/X _12689_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12690_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11641_ _11632_/Y _11633_/X _11634_/Y _11635_/X _11640_/X vssd1 vssd1 vccd1 vccd1
+ _11699_/A sky130_fd_sc_hd__o221a_2
XFILLER_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _14633_/CLK _14360_/D vssd1 vssd1 vccd1 vccd1 _14360_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11572_ _14354_/Q vssd1 vssd1 vccd1 vccd1 _11572_/Y sky130_fd_sc_hd__inv_2
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _14573_/CLK _13311_/D vssd1 vssd1 vccd1 vccd1 _13311_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_in[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_10523_ _13623_/Q vssd1 vssd1 vccd1 vccd1 _10523_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14291_ _14291_/CLK _14291_/D vssd1 vssd1 vccd1 vccd1 _14291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13242_ _13368_/CLK _13242_/D vssd1 vssd1 vccd1 vccd1 _13274_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10454_ _11653_/A vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13173_ _12665_/X _13172_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__mux2_1
X_10385_ _13621_/Q vssd1 vssd1 vccd1 vccd1 _10385_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12124_ vssd1 vssd1 vccd1 vccd1 _12124_/HI _12124_/LO sky130_fd_sc_hd__conb_1
XFILLER_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12055_ _09786_/A _12050_/X _09898_/A _12051_/X vssd1 vssd1 vccd1 vccd1 _12055_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater609 _12658_/S vssd1 vssd1 vccd1 vccd1 _12650_/S sky130_fd_sc_hd__buf_8
X_11006_ _13835_/Q vssd1 vssd1 vccd1 vccd1 _11006_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12558_/X _12956_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11908_ _14089_/Q vssd1 vssd1 vccd1 vccd1 _11908_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12533_/X input337/X _12888_/S vssd1 vssd1 vccd1 vccd1 _12888_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14627_ _14627_/CLK _14627_/D vssd1 vssd1 vccd1 vccd1 _14627_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _14126_/Q vssd1 vssd1 vccd1 vccd1 _11839_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14558_ _14637_/CLK _14558_/D vssd1 vssd1 vccd1 vccd1 _14558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13509_ _14110_/CLK _13509_/D vssd1 vssd1 vccd1 vccd1 _13509_/Q sky130_fd_sc_hd__dfxtp_1
X_14489_ _14611_/CLK _14489_/D vssd1 vssd1 vccd1 vccd1 _14489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07030_ _14553_/Q _07025_/X _06738_/X _07027_/X _07028_/X vssd1 vssd1 vccd1 vccd1
+ _14553_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _08981_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_192_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07932_ _14102_/Q _07926_/X _07778_/X _07927_/X _07929_/X vssd1 vssd1 vccd1 vccd1
+ _14102_/D sky130_fd_sc_hd__o221a_1
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07863_ _07863_/A vssd1 vssd1 vccd1 vccd1 _07863_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06814_ _08167_/A vssd1 vssd1 vccd1 vccd1 _06814_/X sky130_fd_sc_hd__buf_2
X_09602_ _09602_/A vssd1 vssd1 vccd1 vccd1 _12794_/S sky130_fd_sc_hd__inv_16
XFILLER_3_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07794_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09533_ _09533_/A _12415_/X vssd1 vssd1 vccd1 vccd1 _09533_/X sky130_fd_sc_hd__and2_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06745_ _08117_/A vssd1 vssd1 vccd1 vccd1 _06745_/X sky130_fd_sc_hd__buf_2
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09464_ _09479_/A vssd1 vssd1 vccd1 vccd1 _09464_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06676_ _06541_/A _06573_/X _06541_/Y _08912_/A vssd1 vssd1 vccd1 vccd1 _06676_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08415_ _08415_/A vssd1 vssd1 vccd1 vccd1 _08415_/X sky130_fd_sc_hd__clkbuf_2
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09395_ _09395_/A _13135_/X vssd1 vssd1 vccd1 vccd1 _13338_/D sky130_fd_sc_hd__and2_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08346_ _08346_/A vssd1 vssd1 vccd1 vccd1 _08346_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08277_ _13935_/Q _08274_/X _08199_/X _08276_/X _08264_/X vssd1 vssd1 vccd1 vccd1
+ _13935_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07228_ _07262_/A vssd1 vssd1 vccd1 vccd1 _07228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07159_ _08989_/C vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _11042_/A vssd1 vssd1 vccd1 vccd1 _11747_/A sky130_fd_sc_hd__buf_2
XFILLER_106_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput470 _10131_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput481 _12114_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput492 _12124_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13860_ _14095_/CLK _13860_/D vssd1 vssd1 vccd1 vccd1 _13860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _12514_/X _12810_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__mux2_1
X_13791_ _14120_/CLK _13791_/D vssd1 vssd1 vccd1 vccd1 _13791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12742_ _09543_/X _12741_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12742_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _09582_/X _12672_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _13926_/Q vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__inv_2
X_14412_ _14529_/CLK _14412_/D vssd1 vssd1 vccd1 vccd1 _14412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11555_ _11550_/Y _11397_/X _11551_/Y _11399_/X _11554_/X vssd1 vssd1 vccd1 vccd1
+ _11590_/A sky130_fd_sc_hd__o221a_2
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _14627_/CLK _14343_/D vssd1 vssd1 vccd1 vccd1 _14343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _11455_/A vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14274_ _14611_/CLK _14274_/D vssd1 vssd1 vccd1 vccd1 _14274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11486_ _13565_/Q _11430_/X _13806_/Q _11431_/X vssd1 vssd1 vccd1 vccd1 _11486_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13225_ _13352_/CLK _13225_/D vssd1 vssd1 vccd1 vccd1 _13257_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10437_ _10696_/A vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _12657_/X input351/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__mux2_1
X_10368_ _14290_/Q vssd1 vssd1 vccd1 vccd1 _10368_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12107_ vssd1 vssd1 vccd1 vccd1 _12107_/HI _12107_/LO sky130_fd_sc_hd__conb_1
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13087_ _12621_/X _13086_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10299_ _14055_/Q vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__inv_2
X_12038_ _09773_/A _12035_/X _09885_/A _12037_/X vssd1 vssd1 vccd1 vccd1 _12038_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_211_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13989_ _14107_/CLK _13989_/D vssd1 vssd1 vccd1 vccd1 _13989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06530_ _06530_/A vssd1 vssd1 vccd1 vccd1 _06530_/X sky130_fd_sc_hd__buf_2
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08200_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09180_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08131_ _14000_/Q _08122_/X _08130_/X _08124_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _14000_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08062_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07013_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07014_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput209 la_oenb[22] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__buf_1
X_08964_ _13589_/Q _08956_/X _08962_/X _08958_/X _08963_/X vssd1 vssd1 vccd1 vccd1
+ _13589_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _14113_/Q _07910_/X _07751_/X _07911_/X _07913_/X vssd1 vssd1 vccd1 vccd1
+ _14113_/D sky130_fd_sc_hd__o221a_1
XPHY_6518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08895_ _08895_/A vssd1 vssd1 vccd1 vccd1 _08895_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07846_ _07856_/A vssd1 vssd1 vccd1 vccd1 _07846_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07777_ _14181_/Q _07770_/X _07776_/X _07772_/X _07768_/X vssd1 vssd1 vccd1 vccd1
+ _14181_/D sky130_fd_sc_hd__o221a_1
XFILLER_77_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06728_ _09336_/A vssd1 vssd1 vccd1 vccd1 _07130_/A sky130_fd_sc_hd__buf_1
XFILLER_92_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09545_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09450_/A _12983_/X vssd1 vssd1 vccd1 vccd1 _13296_/D sky130_fd_sc_hd__and2_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _06536_/A _08933_/A _06536_/Y _06582_/Y vssd1 vssd1 vccd1 vccd1 _06659_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09378_ _09382_/A _12823_/X vssd1 vssd1 vccd1 vccd1 _13352_/D sky130_fd_sc_hd__and2_1
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08329_ _08329_/A vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11340_ _11335_/Y _11199_/X _11336_/Y _11201_/X _11339_/X vssd1 vssd1 vccd1 vccd1
+ _11353_/B sky130_fd_sc_hd__o221a_1
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _13372_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _11271_/A _11271_/B _11271_/C _11271_/D vssd1 vssd1 vccd1 vccd1 _11271_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_4_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13010_ _13009_/X _12584_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _13010_/X sky130_fd_sc_hd__mux2_1
X_10222_ _11675_/A vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10153_ _10153_/A vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10084_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__buf_2
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13912_ _14146_/CLK _13912_/D vssd1 vssd1 vccd1 vccd1 _13912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13843_ _14110_/CLK _13843_/D vssd1 vssd1 vccd1 vccd1 _13843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13774_ _14094_/CLK _13774_/D vssd1 vssd1 vccd1 vccd1 _13774_/Q sky130_fd_sc_hd__dfxtp_1
X_10986_ _13476_/Q vssd1 vssd1 vccd1 vccd1 _10986_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12725_ _09576_/X _12724_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _09813_/X _13348_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__mux2_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11607_ _13529_/Q vssd1 vssd1 vccd1 vccd1 _11607_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12587_ _09932_/Y _13303_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14326_ _14637_/CLK _14326_/D vssd1 vssd1 vccd1 vccd1 _14326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11538_ _14197_/Q vssd1 vssd1 vccd1 vccd1 _11538_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11469_ _13643_/Q vssd1 vssd1 vccd1 vccd1 _11469_/Y sky130_fd_sc_hd__inv_2
X_14257_ _14305_/CLK _14257_/D vssd1 vssd1 vccd1 vccd1 _14257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13208_ _13368_/CLK _13208_/D vssd1 vssd1 vccd1 vccd1 _13208_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14188_ _14188_/CLK _14188_/D vssd1 vssd1 vccd1 vccd1 _14188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _12647_/X _13138_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07700_ _09131_/A _09063_/B _09201_/C _08673_/D vssd1 vssd1 vccd1 vccd1 _11683_/A
+ sky130_fd_sc_hd__or4_4
X_08680_ _13733_/Q _08677_/X _08589_/X _08679_/X _08671_/X vssd1 vssd1 vccd1 vccd1
+ _13733_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07631_ _07952_/A _10162_/A vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__or2_2
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07562_ _07614_/A vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09301_ _13407_/Q _09294_/X _08132_/A _09295_/X _09298_/X vssd1 vssd1 vccd1 vccd1
+ _13407_/D sky130_fd_sc_hd__o221a_1
X_06513_ _12036_/A vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__buf_6
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07493_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07493_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09232_ _13446_/Q _09224_/X _08927_/X _09225_/X _09228_/X vssd1 vssd1 vccd1 vccd1
+ _13446_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09163_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08114_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _13524_/Q _09086_/X _08927_/X _09087_/X _09093_/X vssd1 vssd1 vccd1 vccd1
+ _13524_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08045_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ _13369_/Q _09996_/B vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__nand2_1
XPHY_7016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _13596_/Q _08944_/X _08945_/X _08946_/X _08938_/X vssd1 vssd1 vccd1 vccd1
+ _13596_/D sky130_fd_sc_hd__o221a_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _13625_/Q _08876_/X _08566_/X _08877_/X _08871_/X vssd1 vssd1 vccd1 vccd1
+ _13625_/D sky130_fd_sc_hd__o221a_1
XFILLER_40_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07829_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ _14066_/Q vssd1 vssd1 vccd1 vccd1 _10840_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _13986_/Q vssd1 vssd1 vccd1 vccd1 _10771_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _13189_/X _13190_/X _12510_/S vssd1 vssd1 vccd1 vccd1 _12510_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13490_ _14291_/CLK _13490_/D vssd1 vssd1 vccd1 vccd1 _13490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12441_ _12440_/X _06909_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12372_ _13214_/Q _12371_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11323_ _13764_/Q vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__inv_2
X_14111_ _14114_/CLK _14111_/D vssd1 vssd1 vccd1 vccd1 _14111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14042_ _14119_/CLK _14042_/D vssd1 vssd1 vccd1 vccd1 _14042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11254_ _14620_/Q vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10205_ _11664_/A vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11185_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _12431_/S sky130_fd_sc_hd__or2_1
XFILLER_136_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10067_ _10102_/B _10113_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__or2_1
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13826_ _14100_/CLK _13826_/D vssd1 vssd1 vccd1 vccd1 _13826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13757_ _13877_/CLK _13757_/D vssd1 vssd1 vccd1 vccd1 _13757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10969_ _11441_/A vssd1 vssd1 vccd1 vccd1 _10969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ _09565_/X input334/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13688_ _14139_/CLK _13688_/D vssd1 vssd1 vccd1 vccd1 _13688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12639_ _13341_/Q _12638_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12639_/X sky130_fd_sc_hd__mux2_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14309_ _14495_/CLK _14309_/D vssd1 vssd1 vccd1 vccd1 _14309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09850_ _09850_/A vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08801_ _08801_/A vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09840_/A sky130_fd_sc_hd__or2_1
X_06993_ _14563_/Q vssd1 vssd1 vccd1 vccd1 _06993_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08732_ _13703_/Q _08730_/X _08566_/X _08731_/X _08728_/X vssd1 vssd1 vccd1 vccd1
+ _13703_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08663_ _08663_/A vssd1 vssd1 vccd1 vccd1 _08663_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07614_ _07614_/A vssd1 vssd1 vccd1 vccd1 _07614_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08594_ _13778_/Q _08588_/X _08490_/X _08591_/X _08592_/X vssd1 vssd1 vccd1 vccd1
+ _13778_/D sky130_fd_sc_hd__o221a_1
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07545_ _14294_/Q _07541_/X _07471_/X _07542_/X _07544_/X vssd1 vssd1 vccd1 vccd1
+ _14294_/D sky130_fd_sc_hd__o221a_1
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07476_ _07476_/A vssd1 vssd1 vccd1 vccd1 _07476_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09215_ _09249_/A vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09077_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08028_ _14052_/Q _08025_/X _07809_/X _08027_/X _08017_/X vssd1 vssd1 vccd1 vccd1
+ _14052_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09979_ _09979_/A vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__inv_2
XPHY_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12989_/X _12574_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _13933_/Q vssd1 vssd1 vccd1 vccd1 _11941_/Y sky130_fd_sc_hd__inv_2
XPHY_6178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ _11867_/Y _10150_/A _11868_/Y _10153_/A _11871_/X vssd1 vssd1 vccd1 vccd1
+ _11907_/A sky130_fd_sc_hd__o221a_2
XPHY_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13611_ _14481_/CLK _13611_/D vssd1 vssd1 vccd1 vccd1 _13611_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10823_ _14377_/Q vssd1 vssd1 vccd1 vccd1 _10823_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ _14621_/CLK _14591_/D vssd1 vssd1 vccd1 vccd1 _14591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _14123_/CLK _13542_/D vssd1 vssd1 vccd1 vccd1 _13542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10754_ _10723_/X _10754_/B _10754_/C _10754_/D vssd1 vssd1 vccd1 vccd1 _10755_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_125_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10685_ _10685_/A _10685_/B _10685_/C _10685_/D vssd1 vssd1 vccd1 vccd1 _10685_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13473_ _14146_/CLK _13473_/D vssd1 vssd1 vccd1 vccd1 _13473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12424_ _12423_/X _06881_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12424_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12355_ _12354_/X _13204_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12355_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11306_ _13919_/Q vssd1 vssd1 vccd1 vccd1 _11306_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12286_ _11948_/Y _14557_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12286_/X sky130_fd_sc_hd__mux2_4
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14025_ _14120_/CLK _14025_/D vssd1 vssd1 vccd1 vccd1 _14025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11237_ _14230_/Q _11170_/X _14425_/Q _11171_/X _11236_/X vssd1 vssd1 vccd1 vccd1
+ _11271_/B sky130_fd_sc_hd__a221oi_2
XFILLER_64_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11168_ _11164_/Y _11165_/X _11166_/Y _11167_/X vssd1 vssd1 vccd1 vccd1 _11168_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10119_ _10126_/A _12457_/X vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11099_ _14500_/Q vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__inv_2
XPHY_7380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13809_ _14121_/CLK _13809_/D vssd1 vssd1 vccd1 vccd1 _13809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07330_ _08117_/A vssd1 vssd1 vccd1 vccd1 _07330_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07261_ _14430_/Q _07257_/X _06760_/X _07258_/X _07254_/X vssd1 vssd1 vccd1 vccd1
+ _14430_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09000_ _09036_/A vssd1 vssd1 vccd1 vccd1 _09000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07192_ _14467_/Q _07185_/X _06766_/X _07186_/X _07189_/X vssd1 vssd1 vccd1 vccd1
+ _14467_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _09902_/A _09937_/A vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__or2_4
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09833_ _09833_/A vssd1 vssd1 vccd1 vccd1 _09833_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09764_ _13324_/Q vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__inv_2
XFILLER_41_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06976_ _06976_/A vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__buf_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08715_ _08723_/A vssd1 vssd1 vccd1 vccd1 _08715_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _09687_/X _09694_/X _09687_/X _09694_/X vssd1 vssd1 vccd1 vccd1 _09695_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08646_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08577_ _08981_/A vssd1 vssd1 vccd1 vccd1 _08577_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_148_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _14304_/Q _07524_/X _07365_/X _07525_/X _07527_/X vssd1 vssd1 vccd1 vccd1
+ _14304_/D sky130_fd_sc_hd__o221a_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07459_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07459_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ _11664_/A vssd1 vssd1 vccd1 vccd1 _11430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09129_ _13501_/Q _09067_/A _08985_/X _09069_/A _09125_/X vssd1 vssd1 vccd1 vccd1
+ _13501_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12140_ vssd1 vssd1 vccd1 vccd1 _12140_/HI _12140_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _09812_/A _12035_/A _09923_/A _09607_/A vssd1 vssd1 vccd1 vccd1 _12071_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_137_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _14303_/Q vssd1 vssd1 vccd1 vccd1 _11022_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _12566_/X _12972_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11924_ _13536_/Q vssd1 vssd1 vccd1 vccd1 _11924_/Y sky130_fd_sc_hd__inv_2
XPHY_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _14204_/Q vssd1 vssd1 vccd1 vccd1 _11855_/Y sky130_fd_sc_hd__inv_2
XPHY_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10806_ _14221_/Q _10696_/X _14416_/Q _10697_/X _10805_/X vssd1 vssd1 vccd1 vccd1
+ _10839_/B sky130_fd_sc_hd__a221oi_2
XFILLER_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14574_ _14595_/CLK _14574_/D vssd1 vssd1 vccd1 vccd1 _14574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_202_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _13650_/Q vssd1 vssd1 vccd1 vccd1 _11786_/Y sky130_fd_sc_hd__inv_2
XPHY_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13525_ _14120_/CLK _13525_/D vssd1 vssd1 vccd1 vccd1 _13525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10737_ _11447_/A vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_207_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13456_ _14169_/CLK _13456_/D vssd1 vssd1 vccd1 vccd1 _13456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10668_ _14608_/Q vssd1 vssd1 vccd1 vccd1 _10668_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12407_ _13218_/Q _06626_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12407_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13387_ _14291_/CLK _13387_/D vssd1 vssd1 vccd1 vccd1 _13387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10599_ _14450_/Q vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ _13193_/Q input92/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ _12059_/Y _13370_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__mux2_1
X_14008_ _14095_/CLK _14008_/D vssd1 vssd1 vccd1 vccd1 _14008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06830_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06761_ _14625_/Q _06751_/X _06760_/X _06754_/X _06749_/X vssd1 vssd1 vccd1 vccd1
+ _14625_/D sky130_fd_sc_hd__o221a_1
XFILLER_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08500_ _08552_/A vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09480_ _09480_/A vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__clkbuf_2
X_06692_ _06853_/B _06691_/A _09060_/A _06691_/Y vssd1 vssd1 vccd1 vccd1 _06692_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08431_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08645_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08362_ _13887_/Q _08354_/X _08119_/X _08356_/X _08359_/X vssd1 vssd1 vccd1 vccd1
+ _13887_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07313_ _07710_/A vssd1 vssd1 vccd1 vccd1 _07313_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08293_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07244_ _07262_/A vssd1 vssd1 vccd1 vccd1 _07244_/X sky130_fd_sc_hd__buf_2
XFILLER_203_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07175_ _07218_/A vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09816_ _09816_/A vssd1 vssd1 vccd1 vccd1 _09816_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09747_ _13341_/Q vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__inv_2
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06959_ _06956_/X _12309_/X _06957_/Y _06958_/X vssd1 vssd1 vccd1 vccd1 _06960_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09678_ _09676_/X _09677_/X _09676_/X _09677_/X vssd1 vssd1 vccd1 vccd1 _09678_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08629_ _13759_/Q _08626_/X _08541_/X _08627_/X _08628_/X vssd1 vssd1 vccd1 vccd1
+ _13759_/D sky130_fd_sc_hd__o221a_1
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11636_/Y _11637_/X _11638_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _11640_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11571_ _14510_/Q vssd1 vssd1 vccd1 vccd1 _11571_/Y sky130_fd_sc_hd__inv_2
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13310_ _14573_/CLK _13310_/D vssd1 vssd1 vccd1 vccd1 _13310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10522_ _13662_/Q vssd1 vssd1 vccd1 vccd1 _10522_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14290_ _14325_/CLK _14290_/D vssd1 vssd1 vccd1 vccd1 _14290_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10453_ _13824_/Q vssd1 vssd1 vccd1 vccd1 _10453_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13241_ _13368_/CLK _13241_/D vssd1 vssd1 vccd1 vccd1 _13273_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_109_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10384_ _13660_/Q vssd1 vssd1 vccd1 vccd1 _10384_/Y sky130_fd_sc_hd__inv_2
X_13172_ _12665_/X input347/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12123_ vssd1 vssd1 vccd1 vccd1 _12123_/HI _12123_/LO sky130_fd_sc_hd__conb_1
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12054_ _09785_/A _12050_/X _09897_/A _12051_/X vssd1 vssd1 vccd1 vccd1 _12054_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_81_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ _11003_/Y _10942_/X _11004_/Y _10944_/X vssd1 vssd1 vccd1 vccd1 _11005_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ _12558_/X input336/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12956_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11907_ _11907_/A _11907_/B _11907_/C _11907_/D vssd1 vssd1 vccd1 vccd1 _11907_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12532_/X _12886_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14627_/CLK _14626_/D vssd1 vssd1 vccd1 vccd1 _14626_/Q sky130_fd_sc_hd__dfxtp_1
X_11838_ _13853_/Q vssd1 vssd1 vccd1 vccd1 _11838_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14557_ _14637_/CLK _14557_/D vssd1 vssd1 vccd1 vccd1 _14557_/Q sky130_fd_sc_hd__dfxtp_1
X_11769_ _14319_/Q vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13508_ _14094_/CLK _13508_/D vssd1 vssd1 vccd1 vccd1 _13508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _14527_/CLK _14488_/D vssd1 vssd1 vccd1 vccd1 _14488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13439_ _14146_/CLK _13439_/D vssd1 vssd1 vccd1 vccd1 _13439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _13582_/Q _08969_/X _08979_/X _08971_/X _08975_/X vssd1 vssd1 vccd1 vccd1
+ _13582_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07931_ _14103_/Q _07926_/X _07776_/X _07927_/X _07929_/X vssd1 vssd1 vccd1 vccd1
+ _14103_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07862_ _14140_/Q _07855_/X _07780_/X _07856_/X _07857_/X vssd1 vssd1 vccd1 vccd1
+ _14140_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09601_ _09601_/A vssd1 vssd1 vccd1 vccd1 _09601_/X sky130_fd_sc_hd__buf_2
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06813_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07793_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07839_/A sky130_fd_sc_hd__buf_4
XFILLER_211_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09530_/X _09528_/X _13281_/Q _09531_/X vssd1 vssd1 vccd1 vccd1 _13249_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_1898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06744_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08117_/A sky130_fd_sc_hd__buf_4
XFILLER_97_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _09500_/A vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__buf_6
X_06675_ _06536_/Y _08927_/A _06536_/A _06645_/Y vssd1 vssd1 vccd1 vccd1 _06675_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08414_ _08468_/A vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ _09395_/A _13131_/X vssd1 vssd1 vccd1 vccd1 _13339_/D sky130_fd_sc_hd__and2_1
XFILLER_40_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08345_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08276_ _08276_/A vssd1 vssd1 vccd1 vccd1 _08276_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07227_ _14445_/Q _07164_/A _06845_/X _07166_/A _07222_/X vssd1 vssd1 vccd1 vccd1
+ _14445_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07158_ _08989_/B vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_133_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ _08660_/A _11669_/A vssd1 vssd1 vccd1 vccd1 _07145_/A sky130_fd_sc_hd__or2_2
XFILLER_156_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput460 _12246_/X vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput471 _10133_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__clkbuf_2
Xoutput482 _12115_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput493 _12125_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12810_ _12514_/X _12809_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12810_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13790_ _14120_/CLK _13790_/D vssd1 vssd1 vccd1 vccd1 _13790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12741_ _09543_/X _12740_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12741_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _09582_/X input358/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12672_/X sky130_fd_sc_hd__mux2_1
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14529_/CLK _14411_/D vssd1 vssd1 vccd1 vccd1 _14411_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11618_/Y _11445_/X _11619_/Y _11447_/X _11622_/X vssd1 vssd1 vccd1 vccd1
+ _11630_/C sky130_fd_sc_hd__o221a_1
XFILLER_106_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _14627_/CLK _14342_/D vssd1 vssd1 vccd1 vccd1 _14342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11554_ _11552_/Y _11401_/X _11553_/Y _11403_/X vssd1 vssd1 vccd1 vccd1 _11554_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11455_/A sky130_fd_sc_hd__buf_6
XFILLER_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ _14611_/CLK _14273_/D vssd1 vssd1 vccd1 vccd1 _14273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _11485_/A vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13224_ _13368_/CLK _13224_/D vssd1 vssd1 vccd1 vccd1 _13256_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_139_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10436_ _10423_/Y _10425_/X _10426_/Y _10428_/X _10435_/X vssd1 vssd1 vccd1 vccd1
+ _10519_/A sky130_fd_sc_hd__o221a_2
XFILLER_136_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13155_ _12655_/X _13154_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__mux2_1
X_10367_ _10362_/Y _10214_/X _10363_/Y _10217_/X _10366_/X vssd1 vssd1 vccd1 vccd1
+ _10380_/B sky130_fd_sc_hd__o221a_2
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12106_ vssd1 vssd1 vccd1 vccd1 _12106_/HI _12106_/LO sky130_fd_sc_hd__conb_1
XFILLER_112_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10298_ _10298_/A _10298_/B _10298_/C _10298_/D vssd1 vssd1 vccd1 vccd1 _10298_/Y
+ sky130_fd_sc_hd__nand4_4
X_13086_ _13085_/X _12621_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12037_ _12065_/A vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__buf_2
XFILLER_120_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13988_ _14107_/CLK _13988_/D vssd1 vssd1 vccd1 vccd1 _13988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12939_ _12549_/X _12938_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14609_ _14627_/CLK _14609_/D vssd1 vssd1 vccd1 vccd1 _14609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08130_ _08130_/A vssd1 vssd1 vccd1 vccd1 _08130_/X sky130_fd_sc_hd__buf_4
XFILLER_202_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08061_ _08069_/A vssd1 vssd1 vccd1 vccd1 _08061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07012_ _07070_/A vssd1 vssd1 vccd1 vccd1 _07069_/A sky130_fd_sc_hd__inv_2
XFILLER_161_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08963_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08963_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07914_ _14114_/Q _07910_/X _07749_/X _07911_/X _07913_/X vssd1 vssd1 vccd1 vccd1
+ _14114_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ _08894_/A vssd1 vssd1 vccd1 vccd1 _08894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07845_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07845_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07776_ _08167_/A vssd1 vssd1 vccd1 vccd1 _07776_/X sky130_fd_sc_hd__buf_4
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _09583_/A vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__inv_2
X_06727_ _09535_/A vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__buf_4
XFILLER_38_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09450_/A _12979_/X vssd1 vssd1 vccd1 vccd1 _13297_/D sky130_fd_sc_hd__and2_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06658_ _06656_/Y _06584_/Y _08950_/A _08965_/A vssd1 vssd1 vccd1 vccd1 _06658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__clkbuf_4
X_06589_ input95/X vssd1 vssd1 vccd1 vccd1 _06589_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08328_ _13905_/Q _08326_/X _08175_/X _08327_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _13905_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08259_ _08259_/A vssd1 vssd1 vccd1 vccd1 _08259_/X sky130_fd_sc_hd__buf_4
XFILLER_166_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _11251_/X _11270_/B _11270_/C _11270_/D vssd1 vssd1 vccd1 vccd1 _11271_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _14365_/Q vssd1 vssd1 vccd1 vccd1 _10221_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _11635_/A vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10083_ _10099_/A _10127_/A vssd1 vssd1 vccd1 vccd1 _12488_/S sky130_fd_sc_hd__or2_1
XFILLER_88_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13911_ _14146_/CLK _13911_/D vssd1 vssd1 vccd1 vccd1 _13911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13842_ _13996_/CLK _13842_/D vssd1 vssd1 vccd1 vccd1 _13842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13773_ _14094_/CLK _13773_/D vssd1 vssd1 vccd1 vccd1 _13773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10985_ _11457_/A vssd1 vssd1 vccd1 vccd1 _10985_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12724_ _09576_/X input361/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _13349_/Q _12654_/X _12655_/S vssd1 vssd1 vccd1 vccd1 _12655_/X sky130_fd_sc_hd__mux2_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11606_ _14004_/Q vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ _13304_/Q _12585_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__mux2_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _14325_/CLK _14325_/D vssd1 vssd1 vccd1 vccd1 _14325_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11537_ _13605_/Q vssd1 vssd1 vccd1 vccd1 _11537_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14256_ _14529_/CLK _14256_/D vssd1 vssd1 vccd1 vccd1 _14256_/Q sky130_fd_sc_hd__dfxtp_1
X_11468_ _13682_/Q vssd1 vssd1 vccd1 vccd1 _11468_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13207_ _13368_/CLK _13207_/D vssd1 vssd1 vccd1 vccd1 _13207_/Q sky130_fd_sc_hd__dfxtp_2
X_10419_ _10417_/Y _10248_/X _10418_/Y _10251_/X vssd1 vssd1 vccd1 vccd1 _10419_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14187_ _14188_/CLK _14187_/D vssd1 vssd1 vccd1 vccd1 _14187_/Q sky130_fd_sc_hd__dfxtp_1
X_11399_ _11399_/A vssd1 vssd1 vccd1 vccd1 _11399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13138_ _13137_/X _12647_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13138_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13069_ _12614_/X _13068_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07630_ _08814_/A _08340_/B _08744_/C _07630_/D vssd1 vssd1 vccd1 vccd1 _10162_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07561_ _07561_/A vssd1 vssd1 vccd1 vccd1 _07561_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09300_ _13408_/Q _09294_/X _08130_/A _09295_/X _09298_/X vssd1 vssd1 vccd1 vccd1
+ _13408_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06512_ _06512_/A _12267_/S vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__or2_1
XFILLER_39_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07492_ _07623_/A vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__buf_2
XFILLER_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09231_ _13447_/Q _09224_/X _08925_/X _09225_/X _09228_/X vssd1 vssd1 vccd1 vccd1
+ _13447_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09162_ _13485_/Q _09155_/X _08927_/X _09156_/X _09157_/X vssd1 vssd1 vccd1 vccd1
+ _13485_/D sky130_fd_sc_hd__o221a_1
XFILLER_72_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08113_ _14008_/Q _08109_/X _08110_/X _08112_/X _08106_/X vssd1 vssd1 vccd1 vccd1
+ _14008_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09093_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08044_ _14043_/Q _08036_/X _07728_/X _08038_/X _08042_/X vssd1 vssd1 vccd1 vccd1
+ _14043_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__inv_2
XPHY_7006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08946_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08946_/X sky130_fd_sc_hd__clkbuf_2
XPHY_7039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _08877_/A vssd1 vssd1 vccd1 vccd1 _08877_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _14160_/Q _07819_/X _07728_/X _07821_/X _07822_/X vssd1 vssd1 vccd1 vccd1
+ _14160_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ _08150_/A vssd1 vssd1 vccd1 vccd1 _07759_/X sky130_fd_sc_hd__buf_4
XPHY_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _10768_/Y _10709_/X _10769_/Y _10711_/X vssd1 vssd1 vccd1 vccd1 _10770_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _09432_/A _13051_/X vssd1 vssd1 vccd1 vccd1 _13311_/D sky130_fd_sc_hd__and2_1
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12440_ _12509_/X _06909_/Y _12440_/S vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _13214_/Q _06639_/A _12416_/S vssd1 vssd1 vccd1 vccd1 _12371_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14110_ _14110_/CLK _14110_/D vssd1 vssd1 vccd1 vccd1 _14110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11322_ _13959_/Q vssd1 vssd1 vccd1 vccd1 _11322_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14119_/CLK _14041_/D vssd1 vssd1 vccd1 vccd1 _14041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11253_ _14347_/Q vssd1 vssd1 vccd1 vccd1 _11253_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10204_ _10204_/A vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__inv_2
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11184_ _14112_/Q vssd1 vssd1 vccd1 vccd1 _11184_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10135_ _10137_/A _12436_/X vssd1 vssd1 vccd1 vccd1 _10135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10066_ _12510_/S _10089_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__or2b_1
XFILLER_27_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13825_ _14100_/CLK _13825_/D vssd1 vssd1 vccd1 vccd1 _13825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13756_ _13877_/CLK _13756_/D vssd1 vssd1 vccd1 vccd1 _13756_/Q sky130_fd_sc_hd__dfxtp_1
X_10968_ _14380_/Q vssd1 vssd1 vccd1 vccd1 _10968_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _09563_/X _12706_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13205_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13687_ _14139_/CLK _13687_/D vssd1 vssd1 vccd1 vccd1 _13687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10899_ _10889_/Y _10702_/X _10892_/X _10895_/X _10898_/X vssd1 vssd1 vccd1 vccd1
+ _10921_/C sky130_fd_sc_hd__o2111a_4
XFILLER_31_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12638_ _09831_/Y _13341_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__mux2_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12569_ _09945_/X _13296_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _14495_/CLK _14308_/D vssd1 vssd1 vccd1 vccd1 _14308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14239_ _14633_/CLK _14239_/D vssd1 vssd1 vccd1 vccd1 _14239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08800_ _08800_/A vssd1 vssd1 vccd1 vccd1 _08800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09780_ _09780_/A _09837_/A vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__or2_1
X_06992_ _06992_/A vssd1 vssd1 vccd1 vccd1 _07004_/A sky130_fd_sc_hd__buf_8
XFILLER_45_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08731_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08731_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08662_ _08662_/A vssd1 vssd1 vccd1 vccd1 _08662_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07613_ _07613_/A vssd1 vssd1 vccd1 vccd1 _07613_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_199_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _13779_/Q _08588_/X _08589_/X _08591_/X _08592_/X vssd1 vssd1 vccd1 vccd1
+ _13779_/D sky130_fd_sc_hd__o221a_1
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07544_ _07576_/A vssd1 vssd1 vccd1 vccd1 _07544_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07475_ _14330_/Q _07467_/X _07396_/X _07468_/X _07469_/X vssd1 vssd1 vccd1 vccd1
+ _14330_/D sky130_fd_sc_hd__o221a_1
XFILLER_201_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09214_ _09257_/A vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__buf_6
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09145_ _09188_/A vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__buf_6
XFILLER_120_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09076_ _09119_/A vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08027_ _08027_/A vssd1 vssd1 vccd1 vccd1 _08027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _13360_/Q _09978_/B vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08929_ _08956_/A vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _11935_/Y _10228_/A _11936_/Y _10231_/A _11939_/X vssd1 vssd1 vccd1 vccd1
+ _11947_/C sky130_fd_sc_hd__o221a_1
XPHY_6168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11871_ _11869_/Y _10156_/A _11870_/Y _10159_/A vssd1 vssd1 vccd1 vccd1 _11871_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13610_ _14481_/CLK _13610_/D vssd1 vssd1 vccd1 vccd1 _13610_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10822_ _14611_/Q vssd1 vssd1 vccd1 vccd1 _10822_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14621_/CLK _14590_/D vssd1 vssd1 vccd1 vccd1 _14590_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13541_ _14123_/CLK _13541_/D vssd1 vssd1 vccd1 vccd1 _13541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10753_ _10744_/Y _10745_/X _10746_/Y _10747_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _10754_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _14146_/CLK _13472_/D vssd1 vssd1 vccd1 vccd1 _13472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10684_ _10665_/X _10684_/B _10684_/C _10684_/D vssd1 vssd1 vccd1 vccd1 _10685_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12423_ _12422_/X _06881_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12423_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ _13204_/Q _12353_/X input78/X vssd1 vssd1 vccd1 vccd1 _12354_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _11300_/Y _11209_/X _11301_/Y _11211_/X _11304_/X vssd1 vssd1 vccd1 vccd1
+ _11312_/C sky130_fd_sc_hd__o221a_1
XFILLER_181_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ _11989_/Y _14558_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12285_/X sky130_fd_sc_hd__mux2_4
XFILLER_153_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14024_ _14119_/CLK _14024_/D vssd1 vssd1 vccd1 vccd1 _14024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11236_ _13404_/Q _11042_/X _13716_/Q _11172_/X vssd1 vssd1 vccd1 vccd1 _11236_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11167_ _11403_/A vssd1 vssd1 vccd1 vccd1 _11167_/X sky130_fd_sc_hd__buf_2
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10118_ _10118_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _12455_/S sky130_fd_sc_hd__or2_1
XFILLER_209_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _13209_/Q _11013_/X _14032_/Q _10957_/X _11097_/X vssd1 vssd1 vccd1 vccd1
+ _11098_/X sky130_fd_sc_hd__a221o_4
XPHY_7370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput360 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input360/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10049_ _13352_/Q _13351_/Q _09966_/A vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _14120_/CLK _13808_/D vssd1 vssd1 vccd1 vccd1 _13808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13739_ _14169_/CLK _13739_/D vssd1 vssd1 vccd1 vccd1 _13739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07260_ _14431_/Q _07257_/X _06757_/X _07258_/X _07254_/X vssd1 vssd1 vccd1 vccd1
+ _14431_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07191_ _14468_/Q _07185_/X _06763_/X _07186_/X _07189_/X vssd1 vssd1 vccd1 vccd1
+ _14468_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__or2_1
XFILLER_47_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ _13342_/Q _09830_/Y _09793_/B vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09763_ _13325_/Q vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__inv_2
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06975_ _14568_/Q vssd1 vssd1 vccd1 vccd1 _06975_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08714_ _08722_/A vssd1 vssd1 vccd1 vccd1 _08714_/X sky130_fd_sc_hd__clkbuf_2
X_09694_ _09656_/A _09693_/X _09656_/A _09693_/X vssd1 vssd1 vccd1 vccd1 _09694_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08645_ _08645_/A vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__clkbuf_4
XPHY_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _13784_/Q _08565_/X _08574_/X _08567_/X _08575_/X vssd1 vssd1 vccd1 vccd1
+ _13784_/D sky130_fd_sc_hd__o221a_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07527_/X sky130_fd_sc_hd__buf_2
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ _14340_/Q _07450_/X _07370_/X _07451_/X _07452_/X vssd1 vssd1 vccd1 vccd1
+ _14340_/D sky130_fd_sc_hd__o221a_1
XFILLER_210_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07389_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07389_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09128_ _13502_/Q _09067_/A _08983_/X _09069_/A _09125_/X vssd1 vssd1 vccd1 vccd1
+ _13502_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09059_ _13540_/Q _08993_/A _08985_/X _08995_/A _09054_/X vssd1 vssd1 vccd1 vccd1
+ _13540_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _09808_/A _12064_/X _09919_/A _12065_/X vssd1 vssd1 vccd1 vccd1 _12070_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _11016_/Y _10963_/X _11017_/Y _10965_/X _11020_/X vssd1 vssd1 vccd1 vccd1
+ _11034_/B sky130_fd_sc_hd__o221a_4
XFILLER_137_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12972_ _12566_/X input332/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12972_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11923_ _14011_/Q vssd1 vssd1 vccd1 vccd1 _11923_/Y sky130_fd_sc_hd__inv_2
XPHY_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _13612_/Q vssd1 vssd1 vccd1 vccd1 _11854_/Y sky130_fd_sc_hd__inv_2
XPHY_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _13395_/Q _10804_/X _13707_/Q _10698_/X vssd1 vssd1 vccd1 vccd1 _10805_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _14573_/CLK _14573_/D vssd1 vssd1 vccd1 vccd1 _14573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ _13689_/Q vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__inv_2
XPHY_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13524_ _14120_/CLK _13524_/D vssd1 vssd1 vccd1 vccd1 _13524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10736_ _13588_/Q vssd1 vssd1 vccd1 vccd1 _10736_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13455_ _14178_/CLK _13455_/D vssd1 vssd1 vccd1 vccd1 _13455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10667_ _14335_/Q vssd1 vssd1 vccd1 vccd1 _10667_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12406_ _12405_/X _13219_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13386_ _14325_/CLK _13386_/D vssd1 vssd1 vccd1 vccd1 _13386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10598_ _13468_/Q vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12337_ _12336_/X _13194_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ _12056_/Y _13369_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14007_ _14095_/CLK _14007_/D vssd1 vssd1 vccd1 vccd1 _14007_/Q sky130_fd_sc_hd__dfxtp_1
X_11219_ _11455_/A vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12199_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06760_ _08128_/A vssd1 vssd1 vccd1 vccd1 _06760_/X sky130_fd_sc_hd__buf_2
XFILLER_168_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput190 la_oenb[120] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__buf_1
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06691_ _06691_/A vssd1 vssd1 vccd1 vccd1 _06691_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08430_ _13850_/Q _08425_/X _08217_/X _08427_/X _08421_/X vssd1 vssd1 vccd1 vccd1
+ _13850_/D sky130_fd_sc_hd__o221a_1
XFILLER_97_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08361_ _13888_/Q _08354_/X _08117_/X _08356_/X _08359_/X vssd1 vssd1 vccd1 vccd1
+ _13888_/D sky130_fd_sc_hd__o221a_1
XFILLER_177_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07312_ _14402_/Q _07307_/X _07311_/X _07309_/X _07301_/X vssd1 vssd1 vccd1 vccd1
+ _14402_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _13926_/Q _08284_/X _08119_/X _08286_/X _08288_/X vssd1 vssd1 vccd1 vccd1
+ _13926_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07243_ _14440_/Q _07238_/X _06719_/X _07240_/X _07228_/X vssd1 vssd1 vccd1 vccd1
+ _14440_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07174_ _07209_/A vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_203_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__or2_1
XFILLER_87_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09746_ _13342_/Q vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__inv_2
XFILLER_60_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06958_ _06958_/A vssd1 vssd1 vccd1 vccd1 _06958_/X sky130_fd_sc_hd__buf_1
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09677_ _06881_/Y _09641_/Y _14593_/Q _09641_/A vssd1 vssd1 vccd1 vccd1 _09677_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06889_ _14591_/Q vssd1 vssd1 vccd1 vccd1 _06889_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08637_/A vssd1 vssd1 vccd1 vccd1 _08628_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08559_ _13791_/Q _08552_/X _08558_/X _08554_/X _08550_/X vssd1 vssd1 vccd1 vccd1
+ _13791_/D sky130_fd_sc_hd__o221a_1
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _13219_/Q _11485_/X _14042_/Q _11429_/X _11569_/X vssd1 vssd1 vccd1 vccd1
+ _11570_/X sky130_fd_sc_hd__a221o_4
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _13428_/Q vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13240_ _13368_/CLK _13240_/D vssd1 vssd1 vccd1 vccd1 _13272_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10452_ _10446_/Y _10448_/X _10449_/Y _10451_/X vssd1 vssd1 vccd1 vccd1 _10452_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13171_ _12663_/X _13170_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10383_ _13426_/Q vssd1 vssd1 vccd1 vccd1 _10383_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ vssd1 vssd1 vccd1 vccd1 _12122_/HI _12122_/LO sky130_fd_sc_hd__conb_1
XFILLER_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12053_ _09784_/A _12050_/X _09896_/A _12051_/X vssd1 vssd1 vccd1 vccd1 _12053_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _13874_/Q vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12955_ _12556_/X _12954_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12955_/X sky130_fd_sc_hd__mux2_1
XPHY_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _11887_/X _11906_/B _11906_/C _11906_/D vssd1 vssd1 vccd1 vccd1 _11907_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12532_/X _12885_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__mux2_1
XPHY_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11837_ _11835_/Y _11648_/X _11836_/Y _11650_/X vssd1 vssd1 vccd1 vccd1 _11837_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _14627_/CLK _14625_/D vssd1 vssd1 vccd1 vccd1 _14625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14556_ _14637_/CLK _14556_/D vssd1 vssd1 vccd1 vccd1 _14556_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11768_ _11763_/Y _11669_/X _11764_/Y _11671_/X _11767_/X vssd1 vssd1 vccd1 vccd1
+ _11781_/B sky130_fd_sc_hd__o221a_2
XFILLER_124_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13507_ _14094_/CLK _13507_/D vssd1 vssd1 vccd1 vccd1 _13507_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10719_ _11429_/A vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__clkbuf_2
X_14487_ _14527_/CLK _14487_/D vssd1 vssd1 vccd1 vccd1 _14487_/Q sky130_fd_sc_hd__dfxtp_1
X_11699_ _11699_/A _11699_/B _11699_/C _11699_/D vssd1 vssd1 vccd1 vccd1 _11699_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13438_ _14146_/CLK _13438_/D vssd1 vssd1 vccd1 vccd1 _13438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13369_ _13371_/CLK _13369_/D vssd1 vssd1 vccd1 vccd1 _13369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07930_ _14104_/Q _07926_/X _07774_/X _07927_/X _07929_/X vssd1 vssd1 vccd1 vccd1
+ _14104_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _14141_/Q _07855_/X _07778_/X _07856_/X _07857_/X vssd1 vssd1 vccd1 vccd1
+ _14141_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ _11485_/A vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__buf_4
XFILLER_116_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06812_ _14611_/Q _06805_/X _06810_/X _06811_/X _06803_/X vssd1 vssd1 vccd1 vccd1
+ _14611_/D sky130_fd_sc_hd__o221a_1
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07792_ _08183_/A vssd1 vssd1 vccd1 vccd1 _07792_/X sky130_fd_sc_hd__buf_4
XFILLER_84_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _09545_/A vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06743_ _06743_/A vssd1 vssd1 vccd1 vccd1 _06743_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09462_ _09501_/A vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__inv_2
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06674_ _06672_/X _06673_/X _06672_/X _06673_/X vssd1 vssd1 vccd1 vccd1 _06674_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ _08469_/A vssd1 vssd1 vccd1 vccd1 _08468_/A sky130_fd_sc_hd__inv_2
X_09393_ _09395_/A _13127_/X vssd1 vssd1 vccd1 vccd1 _13340_/D sky130_fd_sc_hd__and2_1
XFILLER_145_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08344_ _08344_/A vssd1 vssd1 vccd1 vccd1 _08344_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08275_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_197_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07226_ _14446_/Q _07164_/A _06843_/B _07166_/A _07222_/X vssd1 vssd1 vccd1 vccd1
+ _14446_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07157_ _07803_/A vssd1 vssd1 vccd1 vccd1 _08744_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07088_ _07484_/A _07878_/B _08584_/C _07630_/D vssd1 vssd1 vccd1 vccd1 _11669_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput450 _12237_/X vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput461 _12247_/X vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput472 _10135_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput483 _12116_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput494 _12126_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _14595_/Q _09728_/X _14595_/Q _09728_/X vssd1 vssd1 vccd1 vccd1 _09729_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12740_ _09543_/X input343/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _09580_/X _12670_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13198_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14410_ _14529_/CLK _14410_/D vssd1 vssd1 vccd1 vccd1 _14410_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11620_/Y _11449_/X _11621_/Y _11451_/X vssd1 vssd1 vccd1 vccd1 _11622_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _14627_/CLK _14341_/D vssd1 vssd1 vccd1 vccd1 _14341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11553_ _13645_/Q vssd1 vssd1 vccd1 vccd1 _11553_/Y sky130_fd_sc_hd__inv_2
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10504_ _13902_/Q vssd1 vssd1 vccd1 vccd1 _10504_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14272_ _14527_/CLK _14272_/D vssd1 vssd1 vccd1 vccd1 _14272_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11484_ _11474_/Y _11412_/X _11477_/X _11480_/X _11483_/X vssd1 vssd1 vccd1 vccd1
+ _11507_/C sky130_fd_sc_hd__o2111a_4
XFILLER_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13223_ _13368_/CLK _13223_/D vssd1 vssd1 vccd1 vccd1 _13255_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10435_ _10429_/Y _10431_/X _10432_/Y _10434_/X vssd1 vssd1 vccd1 vccd1 _10435_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13154_ _13153_/X _12655_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10364_/Y _10220_/X _10365_/Y _10223_/X vssd1 vssd1 vccd1 vccd1 _10366_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12105_ vssd1 vssd1 vccd1 vccd1 _12105_/HI _12105_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13085_ _12621_/X _13084_/X _13085_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10297_ _10278_/X _10297_/B _10297_/C _10297_/D vssd1 vssd1 vccd1 vccd1 _10298_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_3_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12036_ _12036_/A vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__buf_4
XFILLER_120_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13987_ _14107_/CLK _13987_/D vssd1 vssd1 vccd1 vccd1 _13987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12938_ _12937_/X _12549_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12938_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12528_/X _12868_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14608_ _14611_/CLK _14608_/D vssd1 vssd1 vccd1 vccd1 _14608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14539_ _14595_/CLK _14539_/D vssd1 vssd1 vccd1 vccd1 _14539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08060_ _14033_/Q _08053_/X _07755_/X _08054_/X _08058_/X vssd1 vssd1 vccd1 vccd1
+ _14033_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07011_ _08660_/A _10147_/A vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__or2_2
XFILLER_11_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__buf_4
XFILLER_9_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07913_ _07929_/A vssd1 vssd1 vccd1 vccd1 _07913_/X sky130_fd_sc_hd__buf_2
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08893_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08894_/A sky130_fd_sc_hd__clkbuf_2
XPHY_6509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07844_ _14150_/Q _07837_/X _07755_/X _07838_/X _07839_/X vssd1 vssd1 vccd1 vccd1
+ _14150_/D sky130_fd_sc_hd__o221a_1
XPHY_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07775_ _14182_/Q _07770_/X _07774_/X _07772_/X _07768_/X vssd1 vssd1 vccd1 vccd1
+ _14182_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09583_/A vssd1 vssd1 vccd1 vccd1 _09514_/X sky130_fd_sc_hd__clkbuf_2
X_06726_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06726_/X sky130_fd_sc_hd__buf_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _09445_/A vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__clkbuf_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06657_ _06657_/A vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09376_ _09376_/A _12819_/X vssd1 vssd1 vccd1 vccd1 _13353_/D sky130_fd_sc_hd__and2_1
XFILLER_71_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06588_ input97/X vssd1 vssd1 vccd1 vccd1 _06588_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08327_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08258_ _13944_/Q _08255_/X _08175_/X _08256_/X _08257_/X vssd1 vssd1 vccd1 vccd1
+ _13944_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07209_ _07209_/A vssd1 vssd1 vccd1 vccd1 _07209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08189_ _13977_/Q _08095_/A _08188_/X _08097_/A _08184_/X vssd1 vssd1 vccd1 vccd1
+ _13977_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10220_ _10220_/A vssd1 vssd1 vccd1 vccd1 _10220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10151_ _13422_/Q vssd1 vssd1 vccd1 vccd1 _10151_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10082_ _10107_/B _10122_/A vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__or2_1
XFILLER_87_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13910_ _14143_/CLK _13910_/D vssd1 vssd1 vccd1 vccd1 _13910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13841_ _13996_/CLK _13841_/D vssd1 vssd1 vccd1 vccd1 _13841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13772_ _14094_/CLK _13772_/D vssd1 vssd1 vccd1 vccd1 _13772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _14146_/Q vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12723_ _09573_/X _12722_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13201_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _09817_/Y _13349_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11603_/Y _11419_/X _11604_/Y _11421_/X vssd1 vssd1 vccd1 vccd1 _11605_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _09933_/X _13304_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12585_/X sky130_fd_sc_hd__mux2_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ _14325_/CLK _14324_/D vssd1 vssd1 vccd1 vccd1 _14324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ _14314_/Q vssd1 vssd1 vccd1 vccd1 _11536_/Y sky130_fd_sc_hd__inv_2
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ _14529_/CLK _14255_/D vssd1 vssd1 vccd1 vccd1 _14255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11467_ _13448_/Q vssd1 vssd1 vccd1 vccd1 _11467_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _13368_/CLK _13206_/D vssd1 vssd1 vccd1 vccd1 _13206_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_193_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10418_ _14447_/Q vssd1 vssd1 vccd1 vccd1 _10418_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14186_ _14188_/CLK _14186_/D vssd1 vssd1 vccd1 vccd1 _14186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11398_ _13447_/Q vssd1 vssd1 vccd1 vccd1 _11398_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13137_ _12647_/X _13136_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__mux2_1
X_10349_ _13939_/Q vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13068_ _12614_/X input355/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12019_ _14208_/Q vssd1 vssd1 vccd1 vccd1 _12019_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07560_ _07613_/A vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06511_ _06511_/A vssd1 vssd1 vccd1 vccd1 _12262_/S sky130_fd_sc_hd__buf_6
XFILLER_179_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07491_ _14325_/Q _07488_/X _07412_/X _07490_/X _07476_/X vssd1 vssd1 vccd1 vccd1
+ _14325_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09230_ _13448_/Q _09224_/X _08922_/X _09225_/X _09228_/X vssd1 vssd1 vccd1 vccd1
+ _13448_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _13486_/Q _09155_/X _08925_/X _09156_/X _09157_/X vssd1 vssd1 vccd1 vccd1
+ _13486_/D sky130_fd_sc_hd__o221a_1
XFILLER_206_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08112_ _08163_/A vssd1 vssd1 vccd1 vccd1 _08112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09092_ _09138_/A vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08043_ _14044_/Q _08036_/X _07726_/X _08038_/X _08042_/X vssd1 vssd1 vccd1 vccd1
+ _14044_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _13368_/Q _09994_/B vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ _08945_/A vssd1 vssd1 vccd1 vccd1 _08945_/X sky130_fd_sc_hd__buf_4
XPHY_6306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _08876_/A vssd1 vssd1 vccd1 vccd1 _08876_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _14161_/Q _07819_/X _07726_/X _07821_/X _07822_/X vssd1 vssd1 vccd1 vccd1
+ _14161_/D sky130_fd_sc_hd__o221a_1
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07758_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07758_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06709_ _09535_/A vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07689_ _14217_/Q _07687_/X _07388_/X _07688_/X _07684_/X vssd1 vssd1 vccd1 vccd1
+ _14217_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09428_ _09432_/A _13047_/X vssd1 vssd1 vccd1 vccd1 _13312_/D sky130_fd_sc_hd__and2_1
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09359_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09364_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12370_ _12369_/X _13199_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12370_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _14232_/Q _11170_/X _14427_/Q _11171_/X _11320_/X vssd1 vssd1 vccd1 vccd1
+ _11354_/B sky130_fd_sc_hd__a221oi_2
XFILLER_193_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _14119_/CLK _14040_/D vssd1 vssd1 vccd1 vccd1 _14040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _14503_/Q vssd1 vssd1 vccd1 vccd1 _11252_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _10203_/A vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _11419_/A vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10134_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _12434_/S sky130_fd_sc_hd__or2_1
XFILLER_114_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10065_ _12506_/S _10065_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ _14100_/CLK _13824_/D vssd1 vssd1 vccd1 vccd1 _13824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13755_ _13877_/CLK _13755_/D vssd1 vssd1 vccd1 vccd1 _13755_/Q sky130_fd_sc_hd__dfxtp_1
X_10967_ _11439_/A vssd1 vssd1 vccd1 vccd1 _10967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _09563_/X _12705_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13686_ _14139_/CLK _13686_/D vssd1 vssd1 vccd1 vccd1 _13686_/Q sky130_fd_sc_hd__dfxtp_1
X_10898_ _10896_/Y _10714_/X _10897_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _10898_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_182_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _13342_/Q _12636_/X _12659_/S vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ _13297_/Q _12567_/X input39/X vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _13885_/Q vssd1 vssd1 vccd1 vccd1 _11519_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14307_ _14495_/CLK _14307_/D vssd1 vssd1 vccd1 vccd1 _14307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12499_ _12498_/X _06985_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12499_/X sky130_fd_sc_hd__mux2_2
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14238_ _14633_/CLK _14238_/D vssd1 vssd1 vccd1 vccd1 _14238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14169_ _14169_/CLK _14169_/D vssd1 vssd1 vccd1 vccd1 _14169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06991_ _06991_/A _06991_/B vssd1 vssd1 vccd1 vccd1 _14564_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08730_ _08730_/A vssd1 vssd1 vccd1 vccd1 _08730_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08661_ _08663_/A vssd1 vssd1 vccd1 vccd1 _08662_/A sky130_fd_sc_hd__inv_2
XFILLER_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07612_ _14257_/Q _07605_/X _07383_/X _07606_/X _07609_/X vssd1 vssd1 vccd1 vccd1
+ _14257_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08592_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08592_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07543_ _14295_/Q _07541_/X _07388_/X _07542_/X _07536_/X vssd1 vssd1 vccd1 vccd1
+ _14295_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07474_ _14331_/Q _07467_/X _07394_/X _07468_/X _07469_/X vssd1 vssd1 vccd1 vccd1
+ _14331_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09213_ _13456_/Q _09205_/X _07714_/A _09207_/X _09209_/X vssd1 vssd1 vccd1 vccd1
+ _13456_/D sky130_fd_sc_hd__o221a_1
XFILLER_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09144_ _13495_/Q _09135_/X _08829_/X _09137_/X _09139_/X vssd1 vssd1 vccd1 vccd1
+ _13495_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _13534_/Q _09067_/X _08829_/X _09069_/X _09074_/X vssd1 vssd1 vccd1 vccd1
+ _13534_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08026_ _08079_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09977_ _09977_/A vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__inv_2
XFILLER_58_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _13602_/Q _08916_/X _08927_/X _08918_/X _08923_/X vssd1 vssd1 vccd1 vccd1
+ _13602_/D sky130_fd_sc_hd__o221a_1
XPHY_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08859_ _13636_/Q _08852_/X _08536_/X _08853_/X _08855_/X vssd1 vssd1 vccd1 vccd1
+ _13636_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _13652_/Q vssd1 vssd1 vccd1 vccd1 _11870_/Y sky130_fd_sc_hd__inv_2
XPHY_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10821_ _14338_/Q vssd1 vssd1 vccd1 vccd1 _10821_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13540_ _14123_/CLK _13540_/D vssd1 vssd1 vccd1 vccd1 _13540_/Q sky130_fd_sc_hd__dfxtp_1
X_10752_ _10748_/Y _10749_/X _10750_/Y _10751_/X vssd1 vssd1 vccd1 vccd1 _10752_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _14146_/CLK _13471_/D vssd1 vssd1 vccd1 vccd1 _13471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10683_ _10678_/Y _10506_/X _10679_/Y _10509_/X _10682_/X vssd1 vssd1 vccd1 vccd1
+ _10684_/D sky130_fd_sc_hd__o221a_1
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12422_ _12509_/X _06881_/Y _12422_/S vssd1 vssd1 vccd1 vccd1 _12422_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12353_ _13204_/Q _06603_/A _12368_/S vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ _11302_/Y _11213_/X _11303_/Y _11215_/X vssd1 vssd1 vccd1 vccd1 _11304_/X
+ sky130_fd_sc_hd__o22a_1
X_12284_ _12030_/Y _14559_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12284_/X sky130_fd_sc_hd__mux2_4
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ _14119_/CLK _14023_/D vssd1 vssd1 vccd1 vccd1 _14023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11235_ _11230_/Y _11161_/X _11231_/Y _11163_/X _11234_/X vssd1 vssd1 vccd1 vccd1
+ _11271_/A sky130_fd_sc_hd__o221a_2
XFILLER_153_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11166_ _13637_/Q vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10117_ _10126_/A _12460_/X vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__nor2_8
XFILLER_27_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11097_ _13557_/Q _10958_/X _13798_/Q _10959_/X vssd1 vssd1 vccd1 vccd1 _11097_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_7360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput350 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 input350/X sky130_fd_sc_hd__buf_6
XFILLER_209_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput361 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input361/X sky130_fd_sc_hd__clkbuf_4
XPHY_7382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10048_ _10146_/A _13351_/Q _10116_/A _13351_/Q vssd1 vssd1 vccd1 vccd1 _10048_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13807_ _14120_/CLK _13807_/D vssd1 vssd1 vccd1 vccd1 _13807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _13779_/Q vssd1 vssd1 vccd1 vccd1 _11999_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13738_ _14169_/CLK _13738_/D vssd1 vssd1 vccd1 vccd1 _13738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13669_ _14119_/CLK _13669_/D vssd1 vssd1 vccd1 vccd1 _13669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07190_ _14469_/Q _07185_/X _06760_/X _07186_/X _07189_/X vssd1 vssd1 vccd1 vccd1
+ _14469_/D sky130_fd_sc_hd__o221a_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09900_ _09900_/A _09934_/A vssd1 vssd1 vccd1 vccd1 _09901_/B sky130_fd_sc_hd__or2_1
XFILLER_99_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ _09791_/A _09791_/B _09830_/Y vssd1 vssd1 vccd1 vccd1 _09831_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09762_ _13326_/Q vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__inv_2
X_06974_ _09650_/A vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__buf_1
XFILLER_45_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08713_ _13714_/Q _08706_/X _08536_/X _08707_/X _08712_/X vssd1 vssd1 vccd1 vccd1
+ _13714_/D sky130_fd_sc_hd__o221a_1
X_09693_ _09689_/X _09692_/X _09689_/X _09692_/X vssd1 vssd1 vccd1 vccd1 _09693_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08644_ _08644_/A vssd1 vssd1 vccd1 vccd1 _08644_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08575_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08575_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ _14305_/Q _07524_/X _07362_/X _07525_/X _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14305_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _14341_/Q _07450_/X _07456_/X _07451_/X _07452_/X vssd1 vssd1 vccd1 vccd1
+ _14341_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07388_ _08175_/A vssd1 vssd1 vccd1 vccd1 _07388_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _13503_/Q _09067_/A _08981_/X _09069_/A _09125_/X vssd1 vssd1 vccd1 vccd1
+ _13503_/D sky130_fd_sc_hd__o221a_1
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09058_ _13541_/Q _08993_/A _08983_/X _08995_/A _09054_/X vssd1 vssd1 vccd1 vccd1
+ _13541_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08009_ _14061_/Q _08007_/X _07784_/X _08008_/X _08003_/X vssd1 vssd1 vccd1 vccd1
+ _14061_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11020_ _11018_/Y _10967_/X _11019_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12971_ _12564_/X _12970_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12971_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11920_/Y _10188_/A _11921_/Y _10191_/A vssd1 vssd1 vccd1 vccd1 _11922_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _14321_/Q vssd1 vssd1 vccd1 vccd1 _11853_/Y sky130_fd_sc_hd__inv_2
XPHY_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _11042_/A vssd1 vssd1 vccd1 vccd1 _10804_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11784_ _13455_/Q vssd1 vssd1 vccd1 vccd1 _11784_/Y sky130_fd_sc_hd__inv_2
XPHY_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _14573_/CLK _14572_/D vssd1 vssd1 vccd1 vccd1 _14572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13523_ _14114_/CLK _13523_/D vssd1 vssd1 vccd1 vccd1 _13523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10735_ _11445_/A vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13454_ _14178_/CLK _13454_/D vssd1 vssd1 vccd1 vccd1 _13454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10666_ _14491_/Q vssd1 vssd1 vccd1 vccd1 _10666_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12405_ _13219_/Q _12404_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12405_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13385_ _14325_/CLK _13385_/D vssd1 vssd1 vccd1 vccd1 _13385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10597_ _14138_/Q vssd1 vssd1 vccd1 vccd1 _10597_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _13194_/Q _12335_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12336_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12267_ _12055_/Y _13368_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12267_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14006_ _14095_/CLK _14006_/D vssd1 vssd1 vccd1 vccd1 _14006_/Q sky130_fd_sc_hd__dfxtp_1
X_11218_ _13917_/Q vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__inv_2
X_12198_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11149_ _14267_/Q vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 la_oenb[111] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_hd__buf_1
Xinput191 la_oenb[121] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__buf_1
XFILLER_3_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06690_ _06853_/B vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__clkinv_4
XFILLER_209_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08360_ _13889_/Q _08354_/X _08217_/X _08356_/X _08359_/X vssd1 vssd1 vccd1 vccd1
+ _13889_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07311_ _07708_/A vssd1 vssd1 vccd1 vccd1 _07311_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08291_ _13927_/Q _08284_/X _08117_/X _08286_/X _08288_/X vssd1 vssd1 vccd1 vccd1
+ _13927_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_1920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07242_ _14441_/Q _07238_/X _06714_/X _07240_/X _07228_/X vssd1 vssd1 vccd1 vccd1
+ _14441_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07173_ _07217_/A vssd1 vssd1 vccd1 vccd1 _07209_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _13349_/Q vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__inv_2
XFILLER_115_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09745_ _13343_/Q vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__inv_2
XFILLER_80_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ _14573_/Q vssd1 vssd1 vccd1 vccd1 _06957_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09676_ _09672_/X _09675_/X _09672_/X _09675_/X vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06888_ _06899_/A _06888_/B vssd1 vssd1 vccd1 vccd1 _14592_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08627_ _08636_/A vssd1 vssd1 vccd1 vccd1 _08627_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08558_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08558_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07509_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08489_ _13818_/Q _08486_/X _08199_/X _08488_/X _08480_/X vssd1 vssd1 vccd1 vccd1
+ _13818_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10520_ _14059_/Q vssd1 vssd1 vccd1 vccd1 _10520_/Y sky130_fd_sc_hd__inv_2
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10451_ _11416_/A vssd1 vssd1 vccd1 vccd1 _10451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _13169_/X _12663_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10382_ _14057_/Q vssd1 vssd1 vccd1 vccd1 _10382_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ vssd1 vssd1 vccd1 vccd1 _12121_/HI _12121_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12052_ _09783_/A _12050_/X _09895_/A _12051_/X vssd1 vssd1 vccd1 vccd1 _12052_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11003_ _13757_/Q vssd1 vssd1 vccd1 vccd1 _11003_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12954_ _12953_/X _12556_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__mux2_1
XPHY_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11900_/Y _10242_/A _11901_/Y _10245_/A _11904_/X vssd1 vssd1 vccd1 vccd1
+ _11906_/D sky130_fd_sc_hd__o221a_1
XPHY_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12532_/X _12884_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12885_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14627_/CLK _14624_/D vssd1 vssd1 vccd1 vccd1 _14624_/Q sky130_fd_sc_hd__dfxtp_1
X_11836_ _13892_/Q vssd1 vssd1 vccd1 vccd1 _11836_/Y sky130_fd_sc_hd__inv_2
XPHY_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ _14637_/CLK _14555_/D vssd1 vssd1 vccd1 vccd1 _14555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11765_/Y _11673_/X _11766_/Y _11675_/X vssd1 vssd1 vccd1 vccd1 _11767_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13506_ _14094_/CLK _13506_/D vssd1 vssd1 vccd1 vccd1 _13506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10718_ _10701_/Y _10702_/X _10707_/X _10712_/X _10717_/X vssd1 vssd1 vccd1 vccd1
+ _10755_/C sky130_fd_sc_hd__o2111a_4
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14486_ _14633_/CLK _14486_/D vssd1 vssd1 vccd1 vccd1 _14486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11698_ _11667_/X _11698_/B _11698_/C _11698_/D vssd1 vssd1 vccd1 vccd1 _11699_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_174_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13437_ _14146_/CLK _13437_/D vssd1 vssd1 vccd1 vccd1 _13437_/Q sky130_fd_sc_hd__dfxtp_1
X_10649_ _10647_/Y _10431_/X _10648_/Y _10434_/X vssd1 vssd1 vccd1 vccd1 _10649_/X
+ sky130_fd_sc_hd__o22a_1
X_13368_ _13368_/CLK _13368_/D vssd1 vssd1 vccd1 vccd1 _13368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12319_ _10381_/Y _14524_/Q _12322_/S vssd1 vssd1 vccd1 vccd1 _12319_/X sky130_fd_sc_hd__mux2_4
XFILLER_142_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13299_ _13352_/CLK _13299_/D vssd1 vssd1 vccd1 vccd1 _13299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _14142_/Q _07855_/X _07776_/X _07856_/X _07857_/X vssd1 vssd1 vccd1 vccd1
+ _14142_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06811_ _06811_/A vssd1 vssd1 vccd1 vccd1 _06811_/X sky130_fd_sc_hd__buf_2
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07791_ _14175_/Q _07783_/X _07790_/X _07785_/X _07781_/X vssd1 vssd1 vccd1 vccd1
+ _14175_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06742_ _14630_/Q _06733_/X _06532_/X _08217_/A _06730_/X vssd1 vssd1 vccd1 vccd1
+ _14630_/D sky130_fd_sc_hd__o221a_1
XFILLER_114_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09530_ _09557_/A vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ _13113_/S _09459_/Y _12209_/A _09460_/X vssd1 vssd1 vccd1 vccd1 _09501_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_184_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06673_ _08967_/A _08977_/A _06588_/Y _06574_/Y vssd1 vssd1 vccd1 vccd1 _06673_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08412_ _08745_/A _11653_/A vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__or2_4
X_09392_ _09395_/A _13123_/X vssd1 vssd1 vccd1 vccd1 _13341_/D sky130_fd_sc_hd__and2_1
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ _08396_/A vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08274_ _08274_/A vssd1 vssd1 vccd1 vccd1 _08274_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _14447_/Q _07217_/X _06837_/X _07218_/X _07222_/X vssd1 vssd1 vccd1 vccd1
+ _14447_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07156_ _14482_/Q _07092_/A _07083_/X _07094_/A _07153_/X vssd1 vssd1 vccd1 vccd1
+ _14482_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07087_ _09201_/C vssd1 vssd1 vccd1 vccd1 _08584_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_161_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput440 _12082_/LO vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput451 _12238_/X vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__clkbuf_2
Xoutput462 _12248_/X vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput473 _10137_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__clkbuf_2
Xoutput484 _12117_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_138_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput495 _12127_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07989_ _14073_/Q _07982_/X _07753_/X _07983_/X _07987_/X vssd1 vssd1 vccd1 vccd1
+ _14073_/D sky130_fd_sc_hd__o221a_1
XFILLER_86_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _06886_/Y _14591_/Q _14592_/Q _06889_/Y vssd1 vssd1 vccd1 vccd1 _09728_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09659_ _09657_/X _09658_/X _09657_/X _09658_/X vssd1 vssd1 vccd1 vccd1 _09659_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_186_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _09580_/X _12669_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__mux2_1
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _14277_/Q vssd1 vssd1 vccd1 vccd1 _11621_/Y sky130_fd_sc_hd__inv_2
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _14627_/CLK _14340_/D vssd1 vssd1 vccd1 vccd1 _14340_/Q sky130_fd_sc_hd__dfxtp_1
X_11552_ _13684_/Q vssd1 vssd1 vccd1 vccd1 _11552_/Y sky130_fd_sc_hd__inv_2
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _10490_/Y _10492_/X _10493_/Y _10495_/X _10502_/X vssd1 vssd1 vccd1 vccd1
+ _10518_/C sky130_fd_sc_hd__o221a_1
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11483_ _11481_/Y _11424_/X _11482_/Y _11426_/X vssd1 vssd1 vccd1 vccd1 _11483_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14271_ _14495_/CLK _14271_/D vssd1 vssd1 vccd1 vccd1 _14271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10434_ _11403_/A vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13222_ _13368_/CLK _13222_/D vssd1 vssd1 vccd1 vccd1 _13222_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_193_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10365_ _14368_/Q vssd1 vssd1 vccd1 vccd1 _10365_/Y sky130_fd_sc_hd__inv_2
X_13153_ _12655_/X _13152_/X _13157_/S vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12104_ vssd1 vssd1 vccd1 vccd1 _12104_/HI _12104_/LO sky130_fd_sc_hd__conb_1
XFILLER_65_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13084_ _12621_/X input336/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ _10291_/Y _10242_/X _10292_/Y _10245_/X _10295_/X vssd1 vssd1 vccd1 vccd1
+ _10297_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12035_ _12035_/A vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__buf_2
XFILLER_117_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13986_ _14107_/CLK _13986_/D vssd1 vssd1 vccd1 vccd1 _13986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12937_ _12549_/X _12936_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12528_/X input343/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14629_/CLK _14607_/D vssd1 vssd1 vccd1 vccd1 _14607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11819_ _14476_/Q vssd1 vssd1 vccd1 vccd1 _11819_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ _12511_/X _12798_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12799_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14538_ _14538_/CLK _14538_/D vssd1 vssd1 vccd1 vccd1 _14538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14469_ _14611_/CLK _14469_/D vssd1 vssd1 vccd1 vccd1 _14469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07010_ _07484_/A _07878_/B _08814_/C _07630_/D vssd1 vssd1 vccd1 vccd1 _10147_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _13590_/Q _08956_/X _08960_/X _08958_/X _08951_/X vssd1 vssd1 vccd1 vccd1
+ _13590_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ _14115_/Q _07910_/X _07746_/X _07911_/X _07905_/X vssd1 vssd1 vccd1 vccd1
+ _14115_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08892_ _08971_/A vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__inv_2
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07843_ _14151_/Q _07837_/X _07753_/X _07838_/X _07839_/X vssd1 vssd1 vccd1 vccd1
+ _14151_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07774_ _08165_/A vssd1 vssd1 vccd1 vccd1 _07774_/X sky130_fd_sc_hd__buf_4
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _09847_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09583_/A sky130_fd_sc_hd__or2_4
XFILLER_37_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06725_ _07714_/A vssd1 vssd1 vccd1 vccd1 _06725_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09444_ _09444_/A _12975_/X vssd1 vssd1 vccd1 vccd1 _13298_/D sky130_fd_sc_hd__and2_1
X_06656_ _06657_/A vssd1 vssd1 vccd1 vccd1 _06656_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06587_ _06581_/X _06586_/Y _06581_/X _06586_/Y vssd1 vssd1 vccd1 vccd1 _06587_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09375_ _09376_/A _12815_/X vssd1 vssd1 vccd1 vccd1 _13354_/D sky130_fd_sc_hd__and2_1
XFILLER_178_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08326_ _08326_/A vssd1 vssd1 vccd1 vccd1 _08326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08257_ _08288_/A vssd1 vssd1 vccd1 vccd1 _08257_/X sky130_fd_sc_hd__buf_1
XFILLER_193_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07208_ _14457_/Q _07201_/X _06801_/X _07202_/X _07205_/X vssd1 vssd1 vccd1 vccd1
+ _14457_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _08188_/A vssd1 vssd1 vccd1 vccd1 _08188_/X sky130_fd_sc_hd__buf_4
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07139_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10150_ _10150_/A vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10081_ _10081_/A vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__buf_1
XFILLER_62_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13840_ _13996_/CLK _13840_/D vssd1 vssd1 vccd1 vccd1 _13840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13771_ _14094_/CLK _13771_/D vssd1 vssd1 vccd1 vccd1 _13771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10983_ _11455_/A vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12722_ _09573_/X _12721_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _13350_/Q _12652_/X _12655_/S vssd1 vssd1 vccd1 vccd1 _12653_/X sky130_fd_sc_hd__mux2_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _14121_/Q vssd1 vssd1 vccd1 vccd1 _11604_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _13305_/Q _12583_/X _12647_/S vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__mux2_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _14325_/CLK _14323_/D vssd1 vssd1 vccd1 vccd1 _14323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11535_ _11530_/Y _11435_/X _11531_/Y _11437_/X _11534_/X vssd1 vssd1 vccd1 vccd1
+ _11548_/B sky130_fd_sc_hd__o221a_2
XFILLER_106_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14529_/CLK _14254_/D vssd1 vssd1 vccd1 vccd1 _14254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ _14079_/Q vssd1 vssd1 vccd1 vccd1 _11466_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ _13368_/CLK _13205_/D vssd1 vssd1 vccd1 vccd1 _13205_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_197_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10417_ _13465_/Q vssd1 vssd1 vccd1 vccd1 _10417_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11397_ _11397_/A vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__clkbuf_2
X_14185_ _14305_/CLK _14185_/D vssd1 vssd1 vccd1 vccd1 _14185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _12647_/X input339/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13136_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10348_ _14212_/Q _10164_/X _14407_/Q _10167_/X _10347_/X vssd1 vssd1 vccd1 vccd1
+ _10381_/B sky130_fd_sc_hd__a221oi_2
XFILLER_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10279_ _14483_/Q vssd1 vssd1 vccd1 vccd1 _10279_/Y sky130_fd_sc_hd__inv_2
X_13067_ _12612_/X _13066_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12018_ _13616_/Q vssd1 vssd1 vccd1 vccd1 _12018_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13969_ _14094_/CLK _13969_/D vssd1 vssd1 vccd1 vccd1 _13969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06510_ _06510_/A _09511_/A _06500_/A vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__or3b_1
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07490_ _07490_/A vssd1 vssd1 vccd1 vccd1 _07490_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09160_ _13487_/Q _09155_/X _08922_/X _09156_/X _09157_/X vssd1 vssd1 vccd1 vccd1
+ _13487_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08111_ _08176_/A vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09091_ _13525_/Q _09086_/X _08925_/X _09087_/X _09084_/X vssd1 vssd1 vccd1 vccd1
+ _13525_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08042_ _08066_/A vssd1 vssd1 vccd1 vccd1 _08042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09993_ _09993_/A vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__inv_2
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08944_ _08956_/A vssd1 vssd1 vccd1 vccd1 _08944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08875_ _13626_/Q _08868_/X _08562_/X _08869_/X _08871_/X vssd1 vssd1 vccd1 vccd1
+ _13626_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ _14162_/Q _07819_/X _07825_/X _07821_/X _07822_/X vssd1 vssd1 vccd1 vccd1
+ _14162_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07757_ _14189_/Q _07745_/X _07755_/X _07747_/X _07756_/X vssd1 vssd1 vccd1 vccd1
+ _14189_/D sky130_fd_sc_hd__o221a_1
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06708_ _12282_/X vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__inv_2
X_07688_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07688_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ _09445_/A vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__buf_2
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ _06639_/A vssd1 vssd1 vccd1 vccd1 _06639_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _09509_/A vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__buf_6
XFILLER_16_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08309_ _13916_/Q _08302_/X _08146_/X _08303_/X _08305_/X vssd1 vssd1 vccd1 vccd1
+ _13916_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09289_ _13415_/Q _09285_/X _07723_/A _09287_/X _09280_/X vssd1 vssd1 vccd1 vccd1
+ _13415_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11320_ _13406_/Q _11278_/X _13718_/Q _11172_/X vssd1 vssd1 vccd1 vccd1 _11320_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_125_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _13212_/Q _11249_/X _14035_/Q _11193_/X _11250_/X vssd1 vssd1 vccd1 vccd1
+ _11251_/X sky130_fd_sc_hd__a221o_4
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10202_ _11663_/A vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11182_ _13839_/Q vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _10137_/A _12439_/X vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10064_ _10076_/A _12505_/X vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__nor2_8
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13823_ _14100_/CLK _13823_/D vssd1 vssd1 vccd1 vccd1 _13823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13754_ _13996_/CLK _13754_/D vssd1 vssd1 vccd1 vccd1 _13754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ _14614_/Q vssd1 vssd1 vccd1 vccd1 _10966_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12705_ _09563_/X _12704_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12705_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13685_ _14139_/CLK _13685_/D vssd1 vssd1 vccd1 vccd1 _13685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _13514_/Q vssd1 vssd1 vccd1 vccd1 _10897_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12636_ _09832_/X _13342_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__mux2_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12567_ _09947_/Y _13297_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__mux2_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _14495_/CLK _14306_/D vssd1 vssd1 vccd1 vccd1 _14306_/Q sky130_fd_sc_hd__dfxtp_1
X_11518_ _13768_/Q vssd1 vssd1 vccd1 vccd1 _11518_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12498_ _12497_/X _06985_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__mux2_1
X_14237_ _14611_/CLK _14237_/D vssd1 vssd1 vccd1 vccd1 _14237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11449_ _11449_/A vssd1 vssd1 vccd1 vccd1 _11449_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14168_ _14169_/CLK _14168_/D vssd1 vssd1 vccd1 vccd1 _14168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13119_ _12637_/X _13118_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13119_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14099_ _14100_/CLK _14099_/D vssd1 vssd1 vccd1 vccd1 _14099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06990_ _06974_/X _12318_/X _06989_/X _06976_/X vssd1 vssd1 vccd1 vccd1 _06991_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08660_ _08660_/A _09599_/A vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__or2_2
XFILLER_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07611_ _14258_/Q _07605_/X _07381_/X _07606_/X _07609_/X vssd1 vssd1 vccd1 vccd1
+ _14258_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08591_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07542_ _07542_/A vssd1 vssd1 vccd1 vccd1 _07542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ _14332_/Q _07467_/X _07392_/X _07468_/X _07469_/X vssd1 vssd1 vccd1 vccd1
+ _14332_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09212_ _13457_/Q _09205_/X _07712_/A _09207_/X _09209_/X vssd1 vssd1 vccd1 vccd1
+ _13457_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09143_ _13496_/Q _09135_/X _08827_/X _09137_/X _09139_/X vssd1 vssd1 vccd1 vccd1
+ _13496_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09074_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08025_ _08025_/A vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09976_ _13359_/Q _09976_/B vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08927_ _08927_/A vssd1 vssd1 vccd1 vccd1 _08927_/X sky130_fd_sc_hd__buf_4
XPHY_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _13637_/Q _08852_/X _08534_/X _08853_/X _08855_/X vssd1 vssd1 vccd1 vccd1
+ _13637_/D sky130_fd_sc_hd__o221a_1
XPHY_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07809_ _07809_/A vssd1 vssd1 vccd1 vccd1 _07809_/X sky130_fd_sc_hd__clkbuf_4
XPHY_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08789_ _13672_/Q _08783_/X _08546_/X _08784_/X _08786_/X vssd1 vssd1 vccd1 vccd1
+ _13672_/D sky130_fd_sc_hd__o221a_1
XPHY_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _14494_/Q vssd1 vssd1 vccd1 vccd1 _10820_/Y sky130_fd_sc_hd__inv_2
XPHY_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10751_ _11461_/A vssd1 vssd1 vccd1 vccd1 _10751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13470_ _14146_/CLK _13470_/D vssd1 vssd1 vccd1 vccd1 _13470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10682_ _10680_/Y _10512_/X _10681_/Y _10515_/X vssd1 vssd1 vccd1 vccd1 _10682_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12421_ _12420_/X _06875_/Y _12502_/S vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12352_ _12351_/X _13205_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12352_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11303_ _14270_/Q vssd1 vssd1 vccd1 vccd1 _11303_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12283_ input127/X input295/X _12283_/S vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__mux2_8
XFILLER_194_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14022_ _14047_/CLK _14022_/D vssd1 vssd1 vccd1 vccd1 _14022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11234_ _11232_/Y _11165_/X _11233_/Y _11167_/X vssd1 vssd1 vccd1 vccd1 _11234_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_68_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11165_ _11401_/A vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__buf_2
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10116_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ _11086_/Y _10940_/X _11089_/X _11092_/X _11095_/X vssd1 vssd1 vccd1 vccd1
+ _11118_/C sky130_fd_sc_hd__o2111a_4
XPHY_7350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput340 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input340/X sky130_fd_sc_hd__buf_4
XPHY_7361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput351 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 input351/X sky130_fd_sc_hd__buf_6
XFILLER_27_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ _10128_/A vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__buf_2
Xinput362 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13806_ _14120_/CLK _13806_/D vssd1 vssd1 vccd1 vccd1 _13806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11998_ _13974_/Q vssd1 vssd1 vccd1 vccd1 _11998_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13737_ _14169_/CLK _13737_/D vssd1 vssd1 vccd1 vccd1 _13737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10949_ _11421_/A vssd1 vssd1 vccd1 vccd1 _10949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13668_ _14119_/CLK _13668_/D vssd1 vssd1 vccd1 vccd1 _13668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _13319_/Q _09846_/X _12619_/S vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13599_ _14305_/CLK _13599_/D vssd1 vssd1 vccd1 vccd1 _13599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_0 _10422_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09830_ _09830_/A vssd1 vssd1 vccd1 vccd1 _09830_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _13327_/Q vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__inv_2
XFILLER_132_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06973_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06991_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08712_ _08728_/A vssd1 vssd1 vccd1 vccd1 _08712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09692_ _06872_/Y _09691_/A _14595_/Q _09691_/Y vssd1 vssd1 vccd1 vccd1 _09692_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08643_ _08643_/A vssd1 vssd1 vccd1 vccd1 _08643_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _08979_/A vssd1 vssd1 vccd1 vccd1 _08574_/X sky130_fd_sc_hd__clkbuf_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07525_ _07533_/A vssd1 vssd1 vccd1 vccd1 _07525_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07456_ _08243_/A vssd1 vssd1 vccd1 vccd1 _07456_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07387_ _07387_/A vssd1 vssd1 vccd1 vccd1 _07387_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09126_ _13504_/Q _09119_/X _08979_/X _09120_/X _09125_/X vssd1 vssd1 vccd1 vccd1
+ _13504_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ _13542_/Q _08993_/A _08981_/X _08995_/A _09054_/X vssd1 vssd1 vccd1 vccd1
+ _13542_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08008_ _08008_/A vssd1 vssd1 vccd1 vccd1 _08008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _09884_/A _09884_/B _09958_/Y vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12970_ _12969_/X _12564_/X _13018_/S vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11921_ _14128_/Q vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__inv_2
XPHY_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11852_ _11847_/Y _11669_/X _11848_/Y _11671_/X _11851_/X vssd1 vssd1 vccd1 vccd1
+ _11865_/B sky130_fd_sc_hd__o221a_4
XPHY_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10798_/Y _10687_/X _10799_/Y _10689_/X _10802_/X vssd1 vssd1 vccd1 vccd1
+ _10839_/A sky130_fd_sc_hd__o221a_2
XFILLER_14_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14571_ _14573_/CLK _14571_/D vssd1 vssd1 vccd1 vccd1 _14571_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11783_ _14086_/Q vssd1 vssd1 vccd1 vccd1 _11783_/Y sky130_fd_sc_hd__inv_2
XPHY_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13522_ _14114_/CLK _13522_/D vssd1 vssd1 vccd1 vccd1 _13522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10734_ _14297_/Q vssd1 vssd1 vccd1 vccd1 _10734_/Y sky130_fd_sc_hd__inv_2
XPHY_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13453_ _14178_/CLK _13453_/D vssd1 vssd1 vccd1 vccd1 _13453_/Q sky130_fd_sc_hd__dfxtp_1
X_10665_ _13200_/Q _10539_/X _14023_/Q _10469_/X _10664_/X vssd1 vssd1 vccd1 vccd1
+ _10665_/X sky130_fd_sc_hd__a221o_2
XFILLER_122_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _13219_/Q _06553_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12404_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13384_ _14325_/CLK _13384_/D vssd1 vssd1 vccd1 vccd1 _13384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10596_ _13904_/Q vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12335_ _13194_/Q _06843_/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12266_ _12054_/Y _13367_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12266_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14005_ _14100_/CLK _14005_/D vssd1 vssd1 vccd1 vccd1 _14005_/Q sky130_fd_sc_hd__dfxtp_1
X_11217_ _11208_/Y _11209_/X _11210_/Y _11211_/X _11216_/X vssd1 vssd1 vccd1 vccd1
+ _11228_/C sky130_fd_sc_hd__o221a_1
XFILLER_190_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ _14189_/Q vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11079_ _13440_/Q vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__inv_2
XPHY_7180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput170 la_oenb[102] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__buf_1
XPHY_7191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput181 la_oenb[112] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_hd__buf_1
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput192 la_oenb[122] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__buf_1
XFILLER_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07310_ _14403_/Q _07307_/X _07015_/X _07309_/X _07301_/X vssd1 vssd1 vccd1 vccd1
+ _14403_/D sky130_fd_sc_hd__o221a_1
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08290_ _13928_/Q _08284_/X _08217_/X _08286_/X _08288_/X vssd1 vssd1 vccd1 vccd1
+ _13928_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07241_ _14442_/Q _07238_/X _07015_/X _07240_/X _07228_/X vssd1 vssd1 vccd1 vccd1
+ _14442_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07172_ _14477_/Q _07164_/X _06725_/X _07166_/X _07169_/X vssd1 vssd1 vccd1 vccd1
+ _14477_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput600 _13286_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09813_ _13348_/Q _09809_/Y _09815_/B vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09744_ _12650_/S vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__clkinv_16
XFILLER_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06956_ _06956_/A vssd1 vssd1 vccd1 vccd1 _06956_/X sky130_fd_sc_hd__buf_1
XFILLER_95_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09675_ _09673_/X _09674_/X _09673_/X _09674_/X vssd1 vssd1 vccd1 vccd1 _09675_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06887_ _06880_/X _12290_/X _06886_/Y _06883_/X vssd1 vssd1 vccd1 vccd1 _06888_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08626_ _08635_/A vssd1 vssd1 vccd1 vccd1 _08626_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08557_ _13792_/Q _08552_/X _08556_/X _08554_/X _08550_/X vssd1 vssd1 vccd1 vccd1
+ _13792_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07508_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07508_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08488_ _08488_/A vssd1 vssd1 vccd1 vccd1 _08488_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07439_ _14350_/Q _07432_/X _07345_/X _07433_/X _07434_/X vssd1 vssd1 vccd1 vccd1
+ _14350_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10450_ _11650_/A vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09109_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10381_ _10381_/A _10381_/B _10381_/C _10381_/D vssd1 vssd1 vccd1 vccd1 _10381_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_108_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ vssd1 vssd1 vccd1 vccd1 _12120_/HI _12120_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ _12065_/A vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__buf_4
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _13952_/Q vssd1 vssd1 vccd1 vccd1 _11002_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12953_ _12556_/X _12952_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__mux2_1
XPHY_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _11902_/Y _10248_/A _11903_/Y _10251_/A vssd1 vssd1 vccd1 vccd1 _11904_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12532_/X input338/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__mux2_1
XPHY_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14627_/CLK _14623_/D vssd1 vssd1 vccd1 vccd1 _14623_/Q sky130_fd_sc_hd__dfxtp_1
X_11835_ _13775_/Q vssd1 vssd1 vccd1 vccd1 _11835_/Y sky130_fd_sc_hd__inv_2
XPHY_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14633_/CLK _14554_/D vssd1 vssd1 vccd1 vccd1 _14554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11766_ _14397_/Q vssd1 vssd1 vccd1 vccd1 _11766_/Y sky130_fd_sc_hd__inv_2
XPHY_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13505_ _14094_/CLK _13505_/D vssd1 vssd1 vccd1 vccd1 _13505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10717_ _10713_/Y _10714_/X _10715_/Y _10716_/X vssd1 vssd1 vccd1 vccd1 _10717_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _14637_/CLK _14485_/D vssd1 vssd1 vccd1 vccd1 _14485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11697_ _11688_/Y _11689_/X _11690_/Y _11691_/X _11696_/X vssd1 vssd1 vccd1 vccd1
+ _11698_/D sky130_fd_sc_hd__o221a_1
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13436_ _14146_/CLK _13436_/D vssd1 vssd1 vccd1 vccd1 _13436_/Q sky130_fd_sc_hd__dfxtp_1
X_10648_ _13626_/Q vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13367_ _14639_/CLK _13367_/D vssd1 vssd1 vccd1 vccd1 _13367_/Q sky130_fd_sc_hd__dfxtp_1
X_10579_ _13507_/Q vssd1 vssd1 vccd1 vccd1 _10579_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12318_ _10422_/Y _14525_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13298_ _13877_/CLK _13298_/D vssd1 vssd1 vccd1 vccd1 _13298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12249_ _12249_/A vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06810_ _08165_/A vssd1 vssd1 vccd1 vccd1 _06810_/X sky130_fd_sc_hd__buf_2
X_07790_ _08181_/A vssd1 vssd1 vccd1 vccd1 _07790_/X sky130_fd_sc_hd__buf_4
XFILLER_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06741_ _09009_/A vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__buf_4
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09460_ _12262_/S _09603_/A _09512_/A vssd1 vssd1 vccd1 vccd1 _09460_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06672_ _06600_/Y _06671_/X _06600_/Y _06671_/X vssd1 vssd1 vccd1 vccd1 _06672_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ _08411_/A _09201_/B _08814_/C _08584_/D vssd1 vssd1 vccd1 vccd1 _11653_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_18_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ _09395_/A _13119_/X vssd1 vssd1 vccd1 vccd1 _13342_/D sky130_fd_sc_hd__and2_1
XFILLER_209_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__inv_2
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08273_ _08326_/A vssd1 vssd1 vccd1 vccd1 _08274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07224_ _14448_/Q _07217_/X _06834_/X _07218_/X _07222_/X vssd1 vssd1 vccd1 vccd1
+ _14448_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07155_ _14483_/Q _07092_/A _06850_/B _07094_/A _07153_/X vssd1 vssd1 vccd1 vccd1
+ _14483_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07086_ _07232_/A _07086_/B vssd1 vssd1 vccd1 vccd1 _09201_/C sky130_fd_sc_hd__or2_2
XFILLER_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput430 _12245_/A vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__clkbuf_2
Xoutput441 _12083_/LO vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput452 _12239_/X vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput463 _12249_/X vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__clkbuf_2
Xoutput474 _10139_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput485 _12118_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput496 _12128_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07988_ _14074_/Q _07982_/X _07751_/X _07983_/X _07987_/X vssd1 vssd1 vccd1 vccd1
+ _14074_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09727_ _14593_/Q _09673_/X _14593_/Q _09673_/X vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06939_ _06958_/A vssd1 vssd1 vccd1 vccd1 _06939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09658_ _06886_/Y _14560_/Q _14592_/Q _10057_/A vssd1 vssd1 vccd1 vccd1 _09658_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08609_ _13770_/Q _08599_/X _08510_/X _08601_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _13770_/D sky130_fd_sc_hd__o221a_1
XFILLER_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09597_/A _12334_/X vssd1 vssd1 vccd1 vccd1 _09589_/X sky130_fd_sc_hd__and2_1
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11620_ _14199_/Q vssd1 vssd1 vccd1 vccd1 _11620_/Y sky130_fd_sc_hd__inv_2
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11551_ _13450_/Q vssd1 vssd1 vccd1 vccd1 _11551_/Y sky130_fd_sc_hd__inv_2
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ _10496_/Y _10498_/X _10499_/Y _10501_/X vssd1 vssd1 vccd1 vccd1 _10502_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14495_/CLK _14270_/D vssd1 vssd1 vccd1 vccd1 _14270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11482_ _13526_/Q vssd1 vssd1 vccd1 vccd1 _11482_/Y sky130_fd_sc_hd__inv_2
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13221_ _14188_/CLK _13221_/D vssd1 vssd1 vccd1 vccd1 _13221_/Q sky130_fd_sc_hd__dfxtp_4
X_10433_ _11639_/A vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13152_ _12655_/X input353/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13152_/X sky130_fd_sc_hd__mux2_1
X_10364_ _14602_/Q vssd1 vssd1 vccd1 vccd1 _10364_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ vssd1 vssd1 vccd1 vccd1 _12103_/HI _12103_/LO sky130_fd_sc_hd__conb_1
XFILLER_112_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13083_ _12619_/X _13082_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10295_ _10293_/Y _10248_/X _10294_/Y _10251_/X vssd1 vssd1 vccd1 vccd1 _10295_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _09772_/A _13114_/S _09884_/A _12954_/S vssd1 vssd1 vccd1 vccd1 _12034_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_152_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13985_ _14107_/CLK _13985_/D vssd1 vssd1 vccd1 vccd1 _13985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12936_ _12549_/X input356/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12867_ _12527_/X _12866_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12867_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _13494_/Q vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__inv_2
X_14606_ _14629_/CLK _14606_/D vssd1 vssd1 vccd1 vccd1 _14606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12798_ _12511_/X _12797_/X _12858_/S vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14537_ _14573_/CLK _14537_/D vssd1 vssd1 vccd1 vccd1 _14537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11749_ _13415_/Q _11747_/X _13734_/Q _12416_/S _11748_/X vssd1 vssd1 vccd1 vccd1
+ _11782_/B sky130_fd_sc_hd__a221oi_2
XFILLER_105_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14468_ _14611_/CLK _14468_/D vssd1 vssd1 vccd1 vccd1 _14468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13419_ _14173_/CLK _13419_/D vssd1 vssd1 vccd1 vccd1 _13419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14399_ _14633_/CLK _14399_/D vssd1 vssd1 vccd1 vccd1 _14399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08960_/X sky130_fd_sc_hd__buf_4
XFILLER_48_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07911_ _07927_/A vssd1 vssd1 vccd1 vccd1 _07911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08891_ _09132_/A _11681_/A vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__or2_2
XFILLER_116_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07842_ _14152_/Q _07837_/X _07751_/X _07838_/X _07839_/X vssd1 vssd1 vccd1 vccd1
+ _14152_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07773_ _14183_/Q _07770_/X _07771_/X _07772_/X _07768_/X vssd1 vssd1 vccd1 vccd1
+ _14183_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09512_ _09512_/A _09602_/A vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__or2_1
X_06724_ _08829_/A vssd1 vssd1 vccd1 vccd1 _07714_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09444_/A _12971_/X vssd1 vssd1 vccd1 vccd1 _13299_/D sky130_fd_sc_hd__and2_1
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06655_ _06563_/X _06654_/X _06563_/X _06654_/X vssd1 vssd1 vccd1 vccd1 _06655_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_168_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09374_ _09376_/A _12811_/X vssd1 vssd1 vccd1 vccd1 _13355_/D sky130_fd_sc_hd__and2_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06586_ _06586_/A vssd1 vssd1 vccd1 vccd1 _06586_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08325_ _13906_/Q _08318_/X _08171_/X _08319_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _13906_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08256_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08256_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07207_ _14458_/Q _07201_/X _07058_/X _07202_/X _07205_/X vssd1 vssd1 vccd1 vccd1
+ _14458_/D sky130_fd_sc_hd__o221a_1
X_08187_ _13978_/Q _08095_/A _08186_/X _08097_/A _08184_/X vssd1 vssd1 vccd1 vccd1
+ _13978_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07138_ _14495_/Q _07136_/X _06807_/X _07137_/X _07131_/X vssd1 vssd1 vccd1 vccd1
+ _14495_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07069_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10080_/A _12493_/X vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__nor2_8
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ _14121_/CLK _13770_/D vssd1 vssd1 vccd1 vccd1 _13770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10982_ _13912_/Q vssd1 vssd1 vccd1 vccd1 _10982_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12721_ _09573_/X _12720_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _09819_/X _13350_/Q _12658_/S vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__mux2_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _13848_/Q vssd1 vssd1 vccd1 vccd1 _11603_/Y sky130_fd_sc_hd__inv_2
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12583_ _09935_/Y _13305_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux2_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _14325_/CLK _14322_/D vssd1 vssd1 vccd1 vccd1 _14322_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11534_ _11532_/Y _11439_/X _11533_/Y _11441_/X vssd1 vssd1 vccd1 vccd1 _11534_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14253_ _14529_/CLK _14253_/D vssd1 vssd1 vccd1 vccd1 _14253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11465_ _11465_/A _11465_/B _11465_/C _11465_/D vssd1 vssd1 vccd1 vccd1 _11465_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_125_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _13352_/CLK _13204_/D vssd1 vssd1 vccd1 vccd1 _13204_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_183_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10416_ _14135_/Q vssd1 vssd1 vccd1 vccd1 _10416_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14184_ _14188_/CLK _14184_/D vssd1 vssd1 vccd1 vccd1 _14184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11396_ _14078_/Q vssd1 vssd1 vccd1 vccd1 _11396_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13135_ _12645_/X _13134_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__mux2_1
X_10347_ _13386_/Q _10305_/X _13698_/Q _10173_/X vssd1 vssd1 vccd1 vccd1 _10347_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13066_ _13065_/X _12612_/X _13114_/S vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__mux2_1
X_10278_ _13192_/Q _10276_/X _14015_/Q _10203_/X _10277_/X vssd1 vssd1 vccd1 vccd1
+ _10278_/X sky130_fd_sc_hd__a221o_4
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12017_ _14325_/Q vssd1 vssd1 vccd1 vccd1 _12017_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13968_ _14094_/CLK _13968_/D vssd1 vssd1 vccd1 vccd1 _13968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ _12540_/X _12918_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13899_ _14169_/CLK _13899_/D vssd1 vssd1 vccd1 vccd1 _13899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ _08833_/A vssd1 vssd1 vccd1 vccd1 _08110_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09090_ _13526_/Q _09086_/X _08922_/X _09087_/X _09084_/X vssd1 vssd1 vccd1 vccd1
+ _13526_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08041_ _14045_/Q _08036_/X _07825_/X _08038_/X _08032_/X vssd1 vssd1 vccd1 vccd1
+ _14045_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09992_ _13367_/Q _09992_/B vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08943_ _13597_/Q _08929_/X _08942_/X _08931_/X _08938_/X vssd1 vssd1 vccd1 vccd1
+ _13597_/D sky130_fd_sc_hd__o221a_1
XPHY_7009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ _13627_/Q _08868_/X _08560_/X _08869_/X _08871_/X vssd1 vssd1 vccd1 vccd1
+ _13627_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _08217_/A vssd1 vssd1 vccd1 vccd1 _07825_/X sky130_fd_sc_hd__buf_4
XFILLER_22_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07756_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07756_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06707_ _08895_/A vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__buf_4
XFILLER_129_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07687_ _07687_/A vssd1 vssd1 vccd1 vccd1 _07687_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _09426_/A _13043_/X vssd1 vssd1 vccd1 vccd1 _13313_/D sky130_fd_sc_hd__and2_1
XFILLER_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06638_ _06639_/A vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09357_ _09357_/A _12887_/X vssd1 vssd1 vccd1 vccd1 _13368_/D sky130_fd_sc_hd__and2_1
XFILLER_90_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06569_ _08945_/A vssd1 vssd1 vccd1 vccd1 _06569_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08308_ _13917_/Q _08302_/X _08144_/X _08303_/X _08305_/X vssd1 vssd1 vccd1 vccd1
+ _13917_/D sky130_fd_sc_hd__o221a_1
XFILLER_103_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ _13416_/Q _09285_/X _07719_/A _09287_/X _09280_/X vssd1 vssd1 vccd1 vccd1
+ _13416_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08239_ _08239_/A vssd1 vssd1 vccd1 vccd1 _08239_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _13560_/Q _11194_/X _13801_/Q _11195_/X vssd1 vssd1 vccd1 vccd1 _11250_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _10201_/A vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__inv_2
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11181_ _11177_/Y _11178_/X _11179_/Y _11180_/X vssd1 vssd1 vccd1 vccd1 _11181_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _12437_/S sky130_fd_sc_hd__or2_1
XPHY_7510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10063_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__buf_4
XFILLER_0_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13822_ _14095_/CLK _13822_/D vssd1 vssd1 vccd1 vccd1 _13822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13753_ _13996_/CLK _13753_/D vssd1 vssd1 vccd1 vccd1 _13753_/Q sky130_fd_sc_hd__dfxtp_1
X_10965_ _11437_/A vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__buf_2
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ _09563_/X input335/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13684_ _14143_/CLK _13684_/D vssd1 vssd1 vccd1 vccd1 _13684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _13989_/Q vssd1 vssd1 vccd1 vccd1 _10896_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _13327_/Q _12634_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _13298_/Q _12565_/X input39/X vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _13963_/Q vssd1 vssd1 vccd1 vccd1 _11517_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ _14305_/CLK _14305_/D vssd1 vssd1 vccd1 vccd1 _14305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12497_ _12509_/X _06985_/Y _12497_/S vssd1 vssd1 vccd1 vccd1 _12497_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14236_ _14611_/CLK _14236_/D vssd1 vssd1 vccd1 vccd1 _14236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11448_ _14195_/Q vssd1 vssd1 vccd1 vccd1 _11448_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14167_ _14169_/CLK _14167_/D vssd1 vssd1 vccd1 vccd1 _14167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11379_ _14389_/Q vssd1 vssd1 vccd1 vccd1 _11379_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13118_ _13117_/X _12637_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14098_ _14100_/CLK _14098_/D vssd1 vssd1 vccd1 vccd1 _14098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13049_ _12604_/X _13048_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _13049_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07610_ _14259_/Q _07605_/X _07379_/X _07606_/X _07609_/X vssd1 vssd1 vccd1 vccd1
+ _14259_/D sky130_fd_sc_hd__o221a_1
X_08590_ _08644_/A vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07541_ _07541_/A vssd1 vssd1 vccd1 vccd1 _07541_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07472_ _14333_/Q _07467_/X _07471_/X _07468_/X _07469_/X vssd1 vssd1 vccd1 vccd1
+ _14333_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09211_ _13458_/Q _09205_/X _07710_/A _09207_/X _09209_/X vssd1 vssd1 vccd1 vccd1
+ _13458_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ _13497_/Q _09135_/X _08825_/X _09137_/X _09139_/X vssd1 vssd1 vccd1 vccd1
+ _13497_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09073_ _13535_/Q _09067_/X _08827_/X _09069_/X _09061_/X vssd1 vssd1 vccd1 vccd1
+ _13535_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08024_ _08078_/A vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_198_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _09975_/A vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__inv_2
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08926_ _13603_/Q _08916_/X _08925_/X _08918_/X _08923_/X vssd1 vssd1 vccd1 vccd1
+ _13603_/D sky130_fd_sc_hd__o221a_1
XPHY_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ _13638_/Q _08852_/X _08532_/X _08853_/X _08855_/X vssd1 vssd1 vccd1 vccd1
+ _13638_/D sky130_fd_sc_hd__o221a_1
XPHY_6149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ _07808_/A vssd1 vssd1 vccd1 vccd1 _07808_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08788_ _13673_/Q _08783_/X _08544_/X _08784_/X _08786_/X vssd1 vssd1 vccd1 vccd1
+ _13673_/D sky130_fd_sc_hd__o221a_1
XFILLER_166_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _14196_/Q _07732_/X _07738_/X _07734_/X _07730_/X vssd1 vssd1 vccd1 vccd1
+ _14196_/D sky130_fd_sc_hd__o221a_1
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10750_ _14453_/Q vssd1 vssd1 vccd1 vccd1 _10750_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09409_ _09413_/A _13115_/X vssd1 vssd1 vccd1 vccd1 _13327_/D sky130_fd_sc_hd__and2_1
XFILLER_41_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10681_ _14452_/Q vssd1 vssd1 vccd1 vccd1 _10681_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12420_ _12419_/X _06875_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ _13205_/Q _12350_/X _12396_/S vssd1 vssd1 vccd1 vccd1 _12351_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11302_ _14192_/Q vssd1 vssd1 vccd1 vccd1 _11302_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12282_ input128/X input296/X _12282_/S vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__mux2_8
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14021_ _14047_/CLK _14021_/D vssd1 vssd1 vccd1 vccd1 _14021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11233_ _13638_/Q vssd1 vssd1 vccd1 vccd1 _11233_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11164_ _13676_/Q vssd1 vssd1 vccd1 vccd1 _11164_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _10115_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _12458_/S sky130_fd_sc_hd__or2_1
XFILLER_1_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11095_ _11093_/Y _10952_/X _11094_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput330 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input330/X sky130_fd_sc_hd__buf_6
XPHY_7351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput341 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input341/X sky130_fd_sc_hd__buf_4
X_10046_ _10128_/A vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__buf_2
Xinput352 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input352/X sky130_fd_sc_hd__buf_4
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput363 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__clkbuf_1
XPHY_7384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ _14120_/CLK _13805_/D vssd1 vssd1 vccd1 vccd1 _13805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11997_ _13421_/Q _11747_/A _13740_/Q _09601_/A _11996_/X vssd1 vssd1 vccd1 vccd1
+ _12030_/B sky130_fd_sc_hd__a221oi_2
XPHY_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13736_ _14169_/CLK _13736_/D vssd1 vssd1 vccd1 vccd1 _13736_/Q sky130_fd_sc_hd__dfxtp_1
X_10948_ _14107_/Q vssd1 vssd1 vccd1 vccd1 _10948_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13667_ _14119_/CLK _13667_/D vssd1 vssd1 vccd1 vccd1 _13667_/Q sky130_fd_sc_hd__dfxtp_1
X_10879_ _10860_/X _10879_/B _10879_/C _10879_/D vssd1 vssd1 vccd1 vccd1 _10880_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12618_ _13320_/Q _12617_/X _12619_/S vssd1 vssd1 vccd1 vccd1 _12618_/X sky130_fd_sc_hd__mux2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _14305_/CLK _13598_/D vssd1 vssd1 vccd1 vccd1 _13598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12549_ _13291_/Q _12548_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_1 _10644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14219_ _14470_/CLK _14219_/D vssd1 vssd1 vccd1 vccd1 _14219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09760_ _13328_/Q vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__inv_2
XFILLER_45_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06972_ _06972_/A _06972_/B vssd1 vssd1 vccd1 vccd1 _14569_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08711_ _13715_/Q _08706_/X _08534_/X _08707_/X _08704_/X vssd1 vssd1 vccd1 vccd1
+ _13715_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09691_ _09691_/A vssd1 vssd1 vccd1 vccd1 _09691_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08642_ _13750_/Q _08635_/X _08562_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _13750_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08573_ _13785_/Q _08565_/X _08572_/X _08567_/X _08563_/X vssd1 vssd1 vccd1 vccd1
+ _13785_/D sky130_fd_sc_hd__o221a_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07524_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07524_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07455_ _14342_/Q _07450_/X _07367_/X _07451_/X _07452_/X vssd1 vssd1 vccd1 vccd1
+ _14342_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07386_ _14374_/Q _07373_/X _07383_/X _07375_/X _07385_/X vssd1 vssd1 vccd1 vccd1
+ _14374_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09125_ _09125_/A vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__buf_2
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09056_ _13543_/Q _09048_/X _08979_/X _09049_/X _09054_/X vssd1 vssd1 vccd1 vccd1
+ _13543_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ _08007_/A vssd1 vssd1 vccd1 vccd1 _08007_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_1887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09958_ _09958_/A vssd1 vssd1 vccd1 vccd1 _09958_/Y sky130_fd_sc_hd__inv_2
X_08909_ _13610_/Q _08905_/X _08837_/X _08907_/X _08900_/X vssd1 vssd1 vccd1 vccd1
+ _13610_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09889_/A _09889_/B vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__or2_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _13855_/Q vssd1 vssd1 vccd1 vccd1 _11920_/Y sky130_fd_sc_hd__inv_2
XPHY_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11849_/Y _11673_/X _11850_/Y _11675_/X vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10800_/Y _10691_/X _10801_/Y _10693_/X vssd1 vssd1 vccd1 vccd1 _10802_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14573_/CLK _14570_/D vssd1 vssd1 vccd1 vccd1 _14570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _11782_/A _11782_/B _11782_/C _11782_/D vssd1 vssd1 vccd1 vccd1 _11782_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ _10724_/Y _10725_/X _10726_/Y _10727_/X _10732_/X vssd1 vssd1 vccd1 vccd1
+ _10754_/B sky130_fd_sc_hd__o221a_4
X_13521_ _14114_/CLK _13521_/D vssd1 vssd1 vccd1 vccd1 _13521_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _14178_/CLK _13452_/D vssd1 vssd1 vccd1 vccd1 _13452_/Q sky130_fd_sc_hd__dfxtp_1
X_10664_ _13548_/Q _10471_/X _13789_/Q _10473_/X vssd1 vssd1 vccd1 vccd1 _10664_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12403_ _12402_/X _13220_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12403_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13383_ _14173_/CLK _13383_/D vssd1 vssd1 vccd1 vccd1 _13383_/Q sky130_fd_sc_hd__dfxtp_1
X_10595_ _10590_/Y _10492_/X _10591_/Y _10495_/X _10594_/X vssd1 vssd1 vccd1 vccd1
+ _10602_/C sky130_fd_sc_hd__o221a_1
XFILLER_154_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _12333_/X _13195_/Q _12619_/S vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12265_ _12053_/Y _13366_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12265_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14004_ _14094_/CLK _14004_/D vssd1 vssd1 vccd1 vccd1 _14004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11216_ _11212_/Y _11213_/X _11214_/Y _11215_/X vssd1 vssd1 vccd1 vccd1 _11216_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12196_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11147_ _13597_/Q vssd1 vssd1 vccd1 vccd1 _11147_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _14071_/Q vssd1 vssd1 vccd1 vccd1 _11078_/Y sky130_fd_sc_hd__inv_2
XPHY_7170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput160 la_data_in[94] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_1
XFILLER_209_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput171 la_oenb[103] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__buf_1
XFILLER_3_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10029_ _13381_/Q _10026_/B _10028_/Y _13382_/Q _10026_/Y vssd1 vssd1 vccd1 vccd1
+ _10029_/X sky130_fd_sc_hd__a32o_1
Xinput182 la_oenb[113] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_hd__buf_1
XFILLER_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput193 la_oenb[123] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__buf_1
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13719_ _14183_/CLK _13719_/D vssd1 vssd1 vccd1 vccd1 _13719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07240_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07171_ _14478_/Q _07164_/X _06722_/X _07166_/X _07169_/X vssd1 vssd1 vccd1 vccd1
+ _14478_/D sky130_fd_sc_hd__o221a_1
XFILLER_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput601 _13258_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__or2_1
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09743_ _09743_/A vssd1 vssd1 vccd1 vccd1 _12666_/S sky130_fd_sc_hd__clkbuf_4
X_06955_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06972_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09674_ _06996_/Y _06999_/Y _14562_/Q _14561_/Q vssd1 vssd1 vccd1 vccd1 _09674_/X
+ sky130_fd_sc_hd__a22o_1
X_06886_ _14592_/Q vssd1 vssd1 vccd1 vccd1 _06886_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_41_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08625_ _13760_/Q _08618_/X _08536_/X _08619_/X _08620_/X vssd1 vssd1 vccd1 vccd1
+ _13760_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08556_ _08960_/A vssd1 vssd1 vccd1 vccd1 _08556_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07507_ _14316_/Q _07499_/X _07332_/X _07501_/X _07503_/X vssd1 vssd1 vccd1 vccd1
+ _14316_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08487_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ _14351_/Q _07432_/X _07343_/X _07433_/X _07434_/X vssd1 vssd1 vccd1 vccd1
+ _14351_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07369_ _14380_/Q _07361_/X _07058_/X _07363_/X _07359_/X vssd1 vssd1 vccd1 vccd1
+ _14380_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09108_ _13515_/Q _09103_/X _09035_/X _09104_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _13515_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ _10361_/X _10380_/B _10380_/C _10380_/D vssd1 vssd1 vccd1 vccd1 _10381_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_87_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ _09039_/A vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12050_ _12064_/A vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__buf_4
XFILLER_69_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11001_ _14225_/Q _10933_/X _14420_/Q _10935_/X _11000_/X vssd1 vssd1 vccd1 vccd1
+ _11035_/B sky130_fd_sc_hd__a221oi_2
XFILLER_117_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12952_ _12556_/X input330/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__mux2_1
XPHY_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11903_ _14478_/Q vssd1 vssd1 vccd1 vccd1 _11903_/Y sky130_fd_sc_hd__inv_2
XPHY_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12531_/X _12882_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux2_1
XANTENNA_210 _13283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14622_ _14627_/CLK _14622_/D vssd1 vssd1 vccd1 vccd1 _14622_/Q sky130_fd_sc_hd__dfxtp_1
X_11834_ _13970_/Q vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__inv_2
XPHY_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _14631_/Q vssd1 vssd1 vccd1 vccd1 _11765_/Y sky130_fd_sc_hd__inv_2
X_14553_ _14633_/CLK _14553_/D vssd1 vssd1 vccd1 vccd1 _14553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _14094_/CLK _13504_/D vssd1 vssd1 vccd1 vccd1 _13504_/Q sky130_fd_sc_hd__dfxtp_1
X_10716_ _11426_/A vssd1 vssd1 vccd1 vccd1 _10716_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14484_ _14637_/CLK _14484_/D vssd1 vssd1 vccd1 vccd1 _14484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11696_ _11692_/Y _11693_/X _11694_/Y _11695_/X vssd1 vssd1 vccd1 vccd1 _11696_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10647_ _13665_/Q vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__inv_2
X_13435_ _14143_/CLK _13435_/D vssd1 vssd1 vccd1 vccd1 _13435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13366_ _14639_/CLK _13366_/D vssd1 vssd1 vccd1 vccd1 _13366_/Q sky130_fd_sc_hd__dfxtp_2
X_10578_ _13982_/Q vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12317_ _10519_/Y _14526_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__mux2_2
XFILLER_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13297_ _13352_/CLK _13297_/D vssd1 vssd1 vccd1 vccd1 _13297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12248_ _12248_/A vssd1 vssd1 vccd1 vccd1 _12248_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ vssd1 vssd1 vccd1 vccd1 _12179_/HI _12179_/LO sky130_fd_sc_hd__conb_1
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06740_ _06740_/A vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__inv_2
XFILLER_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06671_ _06545_/Y _06535_/Y _06545_/A _06535_/A vssd1 vssd1 vccd1 vccd1 _06671_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08410_ _08482_/B vssd1 vssd1 vccd1 vccd1 _09201_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__buf_2
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08341_ _08341_/A _11650_/A vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__or2_4
XFILLER_177_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08272_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08326_/A sky130_fd_sc_hd__inv_2
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07223_ _14449_/Q _07217_/X _06831_/X _07218_/X _07222_/X vssd1 vssd1 vccd1 vccd1
+ _14449_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07154_ _14484_/Q _07092_/A _06845_/X _07094_/A _07153_/X vssd1 vssd1 vccd1 vccd1
+ _14484_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07085_ input89/X vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__inv_2
XFILLER_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput420 _12236_/A vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput431 _12246_/A vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput442 _12084_/LO vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput453 _12240_/X vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__clkbuf_2
Xoutput464 _10119_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__clkbuf_2
Xoutput475 _10142_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__clkbuf_2
Xoutput486 _12100_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput497 _12101_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07987_ _08017_/A vssd1 vssd1 vccd1 vccd1 _07987_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09726_/A _10140_/A vssd1 vssd1 vccd1 vccd1 _12508_/S sky130_fd_sc_hd__or2_2
X_06938_ _14578_/Q vssd1 vssd1 vccd1 vccd1 _06938_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _09608_/X _09656_/Y _09608_/X _09656_/Y vssd1 vssd1 vccd1 vccd1 _09657_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06869_ _06869_/A vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08608_ _13771_/Q _08599_/X _08508_/X _08601_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _13771_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09588_ _09588_/A vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__buf_1
XFILLER_103_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _13799_/Q _08526_/X _08536_/X _08528_/X _08538_/X vssd1 vssd1 vccd1 vccd1
+ _13799_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _14081_/Q vssd1 vssd1 vccd1 vccd1 _11550_/Y sky130_fd_sc_hd__inv_2
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ _11451_/A vssd1 vssd1 vccd1 vccd1 _10501_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11481_ _14001_/Q vssd1 vssd1 vccd1 vccd1 _11481_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13220_ _13350_/CLK _13220_/D vssd1 vssd1 vccd1 vccd1 _13220_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10432_ _13622_/Q vssd1 vssd1 vccd1 vccd1 _10432_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13151_ _12653_/X _13150_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13151_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _14329_/Q vssd1 vssd1 vccd1 vccd1 _10363_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ vssd1 vssd1 vccd1 vccd1 _12102_/HI _12102_/LO sky130_fd_sc_hd__conb_1
XFILLER_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ _13081_/X _12619_/X _13146_/S vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__mux2_1
X_10294_ _14444_/Q vssd1 vssd1 vccd1 vccd1 _10294_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12033_ _09771_/A _13114_/S _09883_/A _12954_/S vssd1 vssd1 vccd1 vccd1 _12033_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_156_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _14107_/CLK _13984_/D vssd1 vssd1 vccd1 vccd1 _13984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12935_ _12547_/X _12934_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12527_/X _12865_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14605_ _14629_/CLK _14605_/D vssd1 vssd1 vccd1 vccd1 _14605_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11817_ _14164_/Q vssd1 vssd1 vccd1 vccd1 _11817_/Y sky130_fd_sc_hd__inv_2
XPHY_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12797_ _12511_/X _12796_/X _12853_/S vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14536_ _14595_/CLK _14536_/D vssd1 vssd1 vccd1 vccd1 _14536_/Q sky130_fd_sc_hd__dfxtp_1
X_11748_ _14241_/Q _11406_/A _14436_/Q _11407_/A vssd1 vssd1 vccd1 vccd1 _11748_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_174_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14467_ _14611_/CLK _14467_/D vssd1 vssd1 vccd1 vccd1 _14467_/Q sky130_fd_sc_hd__dfxtp_1
X_11679_ _11679_/A vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__buf_2
XFILLER_204_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13418_ _14173_/CLK _13418_/D vssd1 vssd1 vccd1 vccd1 _13418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14398_ _14633_/CLK _14398_/D vssd1 vssd1 vccd1 vccd1 _14398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13349_ _13350_/CLK _13349_/D vssd1 vssd1 vccd1 vccd1 _13349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07910_ _07926_/A vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08890_ _09271_/A _08890_/B _09201_/C _09201_/D vssd1 vssd1 vccd1 vccd1 _11681_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_83_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07841_ _14153_/Q _07837_/X _07749_/X _07838_/X _07839_/X vssd1 vssd1 vccd1 vccd1
+ _14153_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07772_ _07772_/A vssd1 vssd1 vccd1 vccd1 _07772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06723_ _14634_/Q _06530_/X _06722_/X _06716_/X _06723_/C1 vssd1 vssd1 vccd1 vccd1
+ _14634_/D sky130_fd_sc_hd__o221a_1
X_09511_ _09511_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09602_/A sky130_fd_sc_hd__or2_4
XFILLER_42_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09442_ _09444_/A _12967_/X vssd1 vssd1 vccd1 vccd1 _13300_/D sky130_fd_sc_hd__and2_1
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06654_ _08985_/A _06653_/X _06608_/A _06653_/X vssd1 vssd1 vccd1 vccd1 _06654_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09373_ _09376_/A _12807_/X vssd1 vssd1 vccd1 vccd1 _13356_/D sky130_fd_sc_hd__and2_1
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06585_ _06582_/Y _08965_/A _06609_/A _06584_/Y vssd1 vssd1 vccd1 vccd1 _06586_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08324_ _13907_/Q _08318_/X _08169_/X _08319_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _13907_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08255_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08255_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07206_ _14459_/Q _07201_/X _06796_/X _07202_/X _07205_/X vssd1 vssd1 vccd1 vccd1
+ _14459_/D sky130_fd_sc_hd__o221a_1
XFILLER_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08186_ _08186_/A vssd1 vssd1 vccd1 vccd1 _08186_/X sky130_fd_sc_hd__buf_4
XFILLER_140_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07137_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07068_ _14530_/Q _07061_/X _06820_/X _07062_/X _07063_/X vssd1 vssd1 vccd1 vccd1
+ _14530_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _09688_/X _09708_/X _09688_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10981_ _10972_/Y _10973_/X _10974_/Y _10975_/X _10980_/X vssd1 vssd1 vccd1 vccd1
+ _10992_/C sky130_fd_sc_hd__o221a_1
XFILLER_99_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _09573_/X input331/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12720_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _13335_/Q _12650_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11600_/Y _11414_/X _11601_/Y _11416_/X vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12582_ _13306_/Q _12581_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12582_/X sky130_fd_sc_hd__mux2_1
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ _14325_/CLK _14321_/D vssd1 vssd1 vccd1 vccd1 _14321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _14392_/Q vssd1 vssd1 vccd1 vccd1 _11533_/Y sky130_fd_sc_hd__inv_2
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _14291_/CLK _14252_/D vssd1 vssd1 vccd1 vccd1 _14252_/Q sky130_fd_sc_hd__dfxtp_1
X_11464_ _11433_/X _11464_/B _11464_/C _11464_/D vssd1 vssd1 vccd1 vccd1 _11465_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_172_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10415_ _13901_/Q vssd1 vssd1 vccd1 vccd1 _10415_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13203_ _13352_/CLK _13203_/D vssd1 vssd1 vccd1 vccd1 _13203_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_171_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11395_ _11395_/A _11395_/B _11395_/C _11395_/D vssd1 vssd1 vccd1 vccd1 _11395_/Y
+ sky130_fd_sc_hd__nand4_4
X_14183_ _14183_/CLK _14183_/D vssd1 vssd1 vccd1 vccd1 _14183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10341_/Y _10150_/X _10342_/Y _10153_/X _10345_/X vssd1 vssd1 vccd1 vccd1
+ _10381_/A sky130_fd_sc_hd__o221a_2
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13134_ _13133_/X _12645_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13065_ _12612_/X _13064_/X _13109_/S vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10277_ _13540_/Q _10206_/X _13781_/Q _10209_/X vssd1 vssd1 vccd1 vccd1 _10277_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12016_ _12011_/Y _10214_/A _12012_/Y _10217_/A _12015_/X vssd1 vssd1 vccd1 vccd1
+ _12029_/B sky130_fd_sc_hd__o221a_4
XFILLER_191_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13967_ _14094_/CLK _13967_/D vssd1 vssd1 vccd1 vccd1 _13967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _12540_/X _12917_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12918_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13898_ _14169_/CLK _13898_/D vssd1 vssd1 vccd1 vccd1 _13898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ _12523_/X _12848_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14519_ _14637_/CLK _14519_/D vssd1 vssd1 vccd1 vccd1 _14519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08040_ _14046_/Q _08036_/X _07723_/X _08038_/X _08032_/X vssd1 vssd1 vccd1 vccd1
+ _14046_/D sky130_fd_sc_hd__o221a_1
XFILLER_89_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09991_ _09991_/A vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__inv_2
XFILLER_142_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08942_ _08942_/A vssd1 vssd1 vccd1 vccd1 _08942_/X sky130_fd_sc_hd__buf_6
XFILLER_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08873_ _13628_/Q _08868_/X _08558_/X _08869_/X _08871_/X vssd1 vssd1 vccd1 vccd1
+ _13628_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07824_ _14163_/Q _07819_/X _07723_/X _07821_/X _07822_/X vssd1 vssd1 vccd1 vccd1
+ _14163_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07755_ _08146_/A vssd1 vssd1 vccd1 vccd1 _07755_/X sky130_fd_sc_hd__buf_4
XPHY_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06706_ _06743_/A _06705_/X _06743_/A _06705_/X vssd1 vssd1 vccd1 vccd1 _08895_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07686_ _14218_/Q _07679_/X _07383_/X _07680_/X _07684_/X vssd1 vssd1 vccd1 vccd1
+ _14218_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09425_ _09426_/A _13039_/X vssd1 vssd1 vccd1 vccd1 _13314_/D sky130_fd_sc_hd__and2_1
X_06637_ input96/X vssd1 vssd1 vccd1 vccd1 _06637_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09356_ _09357_/A _12883_/X vssd1 vssd1 vccd1 vccd1 _13369_/D sky130_fd_sc_hd__and2_1
X_06568_ _06544_/Y _06696_/A _06546_/A _06567_/Y vssd1 vssd1 vccd1 vccd1 _06568_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08307_ _13918_/Q _08302_/X _08142_/X _08303_/X _08305_/X vssd1 vssd1 vccd1 vccd1
+ _13918_/D sky130_fd_sc_hd__o221a_1
XFILLER_205_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09287_ _09319_/A vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__clkbuf_2
X_06499_ _06499_/A _06499_/B _06499_/C _06499_/D vssd1 vssd1 vccd1 vccd1 _06510_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08238_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08169_ _08169_/A vssd1 vssd1 vccd1 vccd1 _08169_/X sky130_fd_sc_hd__buf_4
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10200_ _10176_/Y _10178_/X _10185_/X _10192_/X _10199_/X vssd1 vssd1 vccd1 vccd1
+ _10255_/C sky130_fd_sc_hd__o2111a_4
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _11416_/A vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10131_ _10137_/A _12442_/X vssd1 vssd1 vccd1 vccd1 _10131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10079_/A _10145_/A vssd1 vssd1 vccd1 vccd1 _12503_/S sky130_fd_sc_hd__or2_1
XPHY_7533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ _14095_/CLK _13821_/D vssd1 vssd1 vccd1 vccd1 _13821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13752_ _13996_/CLK _13752_/D vssd1 vssd1 vccd1 vccd1 _13752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10964_ _14341_/Q vssd1 vssd1 vccd1 vccd1 _10964_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12703_ _09560_/X _12702_/X _13155_/S vssd1 vssd1 vccd1 vccd1 _13206_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13683_ _14143_/CLK _13683_/D vssd1 vssd1 vccd1 vccd1 _13683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10895_ _10893_/Y _10709_/X _10894_/Y _10711_/X vssd1 vssd1 vccd1 vccd1 _10895_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _09834_/Y _13327_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12565_ _09948_/X _13298_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__mux2_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _14305_/CLK _14304_/D vssd1 vssd1 vccd1 vccd1 _14304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11516_ _14236_/Q _11406_/X _14431_/Q _11407_/X _11515_/X vssd1 vssd1 vccd1 vccd1
+ _11549_/B sky130_fd_sc_hd__a221oi_2
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12495_/X _06982_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__mux2_2
XFILLER_201_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14235_ _14611_/CLK _14235_/D vssd1 vssd1 vccd1 vccd1 _14235_/Q sky130_fd_sc_hd__dfxtp_1
X_11447_ _11447_/A vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14166_ _14169_/CLK _14166_/D vssd1 vssd1 vccd1 vccd1 _14166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11378_ _14623_/Q vssd1 vssd1 vccd1 vccd1 _11378_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10329_ _14172_/Q vssd1 vssd1 vccd1 vccd1 _10329_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ _12637_/X _13116_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_14097_ _14100_/CLK _14097_/D vssd1 vssd1 vccd1 vccd1 _14097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13048_ _12604_/X input346/X _13176_/S vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07540_ _14296_/Q _07532_/X _07383_/X _07533_/X _07536_/X vssd1 vssd1 vccd1 vccd1
+ _14296_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07471_ _08259_/A vssd1 vssd1 vccd1 vccd1 _07471_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09210_ _13459_/Q _09205_/X _07708_/A _09207_/X _09209_/X vssd1 vssd1 vccd1 vccd1
+ _13459_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ _13498_/Q _09135_/X _08822_/X _09137_/X _09139_/X vssd1 vssd1 vccd1 vccd1
+ _13498_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09072_ _13536_/Q _09067_/X _08825_/X _09069_/X _09061_/X vssd1 vssd1 vccd1 vccd1
+ _13536_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08023_ _08079_/A vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__inv_2
XFILLER_198_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _13358_/Q _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08925_ _08925_/A vssd1 vssd1 vccd1 vccd1 _08925_/X sky130_fd_sc_hd__buf_6
XFILLER_83_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08856_ _13639_/Q _08852_/X _08530_/X _08853_/X _08855_/X vssd1 vssd1 vccd1 vccd1
+ _13639_/D sky130_fd_sc_hd__o221a_1
XPHY_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07807_ _07863_/A vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__clkbuf_2
XPHY_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08787_ _13674_/Q _08783_/X _08541_/X _08784_/X _08786_/X vssd1 vssd1 vccd1 vccd1
+ _13674_/D sky130_fd_sc_hd__o221a_1
XPHY_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _08128_/A vssd1 vssd1 vccd1 vccd1 _07738_/X sky130_fd_sc_hd__buf_4
XPHY_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07669_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07669_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _09414_/A vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__clkbuf_2
X_10680_ _13470_/Q vssd1 vssd1 vccd1 vccd1 _10680_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09339_ _13383_/Q _09275_/A _09060_/X _09277_/A _09352_/A vssd1 vssd1 vccd1 vccd1
+ _13383_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12350_ _13205_/Q _06558_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11301_ _13600_/Q vssd1 vssd1 vccd1 vccd1 _11301_/Y sky130_fd_sc_hd__inv_2
X_12281_ _12073_/Y _13382_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12281_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14020_ _14047_/CLK _14020_/D vssd1 vssd1 vccd1 vccd1 _14020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11232_ _13677_/Q vssd1 vssd1 vccd1 vccd1 _11232_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11163_ _11399_/A vssd1 vssd1 vccd1 vccd1 _11163_/X sky130_fd_sc_hd__buf_2
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10114_/A _12463_/X vssd1 vssd1 vccd1 vccd1 _12248_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11094_ _13518_/Q vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__inv_2
XPHY_7330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput320 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _06497_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput331 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 input331/X sky130_fd_sc_hd__clkbuf_4
XPHY_7352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10045_ _13366_/Q _09990_/B _09991_/A vssd1 vssd1 vccd1 vccd1 _10045_/X sky130_fd_sc_hd__o21a_1
Xinput342 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input342/X sky130_fd_sc_hd__buf_4
XPHY_7363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput353 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 input353/X sky130_fd_sc_hd__buf_6
XPHY_7374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput364 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__clkbuf_1
XPHY_7385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _14120_/CLK _13804_/D vssd1 vssd1 vccd1 vccd1 _13804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11996_ _14247_/Q _11830_/X _14442_/Q _11831_/X vssd1 vssd1 vccd1 vccd1 _11996_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_166_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13735_ _14169_/CLK _13735_/D vssd1 vssd1 vccd1 vccd1 _13735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _11419_/A vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13666_ _14119_/CLK _13666_/D vssd1 vssd1 vccd1 vccd1 _13666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10878_ _10873_/Y _10745_/X _10874_/Y _10747_/X _10877_/X vssd1 vssd1 vccd1 vccd1
+ _10879_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _09848_/X _13320_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12617_/X sky130_fd_sc_hd__mux2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _14305_/CLK _13597_/D vssd1 vssd1 vccd1 vccd1 _13597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12548_ _09960_/X _13291_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_2 _10685_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12509_/X _06961_/Y _12479_/S vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14218_ _14470_/CLK _14218_/D vssd1 vssd1 vccd1 vccd1 _14218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14149_ _14188_/CLK _14149_/D vssd1 vssd1 vccd1 vccd1 _14149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06971_ _06956_/X _12313_/X _06970_/Y _06958_/X vssd1 vssd1 vccd1 vccd1 _06972_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08710_ _13716_/Q _08706_/X _08532_/X _08707_/X _08704_/X vssd1 vssd1 vccd1 vccd1
+ _13716_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09690_ _06989_/A _14563_/Q _14564_/Q _06993_/Y vssd1 vssd1 vccd1 vccd1 _09691_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08641_ _13751_/Q _08635_/X _08560_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _13751_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08572_ _08977_/A vssd1 vssd1 vccd1 vccd1 _08572_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07523_ _14306_/Q _07516_/X _07358_/X _07517_/X _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14306_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07454_ _14343_/Q _07450_/X _07365_/X _07451_/X _07452_/X vssd1 vssd1 vccd1 vccd1
+ _14343_/D sky130_fd_sc_hd__o221a_1
XFILLER_91_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07385_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07385_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _13505_/Q _09119_/X _08977_/X _09120_/X _09117_/X vssd1 vssd1 vccd1 vccd1
+ _13505_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09055_ _13544_/Q _09048_/X _08977_/X _09049_/X _09054_/X vssd1 vssd1 vccd1 vccd1
+ _13544_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ _14062_/Q _07999_/X _07780_/X _08000_/X _08003_/X vssd1 vssd1 vccd1 vccd1
+ _14062_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09883_/A _09883_/B _09884_/B vssd1 vssd1 vccd1 vccd1 _09957_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08908_ _13611_/Q _08905_/X _08833_/X _08907_/X _08900_/X vssd1 vssd1 vccd1 vccd1
+ _13611_/D sky130_fd_sc_hd__o221a_1
XFILLER_8_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09888_ _09888_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09889_/B sky130_fd_sc_hd__or2_1
XFILLER_150_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08871_/A vssd1 vssd1 vccd1 vccd1 _08839_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11850_ _14399_/Q vssd1 vssd1 vccd1 vccd1 _11850_/Y sky130_fd_sc_hd__inv_2
XPHY_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _13629_/Q vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11781_ _11762_/X _11781_/B _11781_/C _11781_/D vssd1 vssd1 vccd1 vccd1 _11782_/D
+ sky130_fd_sc_hd__and4b_2
XPHY_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _14114_/CLK _13520_/D vssd1 vssd1 vccd1 vccd1 _13520_/Q sky130_fd_sc_hd__dfxtp_1
X_10732_ _10728_/Y _10729_/X _10730_/Y _10731_/X vssd1 vssd1 vccd1 vccd1 _10732_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13451_ _14178_/CLK _13451_/D vssd1 vssd1 vccd1 vccd1 _13451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10663_ _10653_/Y _10445_/X _10656_/X _10659_/X _10662_/X vssd1 vssd1 vccd1 vccd1
+ _10685_/C sky130_fd_sc_hd__o2111a_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12402_ _13220_/Q _12401_/X _12417_/S vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ _10592_/Y _10498_/X _10593_/Y _10501_/X vssd1 vssd1 vccd1 vccd1 _10594_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13382_ _14538_/CLK _13382_/D vssd1 vssd1 vccd1 vccd1 _13382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12333_ _13195_/Q _12332_/X input78/X vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12264_ _12052_/Y _13365_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _14110_/CLK _14003_/D vssd1 vssd1 vccd1 vccd1 _14003_/Q sky130_fd_sc_hd__dfxtp_1
X_11215_ _11451_/A vssd1 vssd1 vccd1 vccd1 _11215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12195_ vssd1 vssd1 vccd1 vccd1 _12195_/HI _12195_/LO sky130_fd_sc_hd__conb_1
XFILLER_64_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11146_ _14306_/Q vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11077_ _11077_/A _11077_/B _11077_/C _11077_/D vssd1 vssd1 vccd1 vccd1 _11077_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_62_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput150 la_data_in[85] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__buf_1
XPHY_7171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput161 la_data_in[95] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_1
XFILLER_23_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10028_ _13382_/Q vssd1 vssd1 vccd1 vccd1 _10028_/Y sky130_fd_sc_hd__inv_2
Xinput172 la_oenb[104] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_hd__buf_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput183 la_oenb[114] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__buf_1
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput194 la_oenb[124] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__buf_1
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11979_ _14285_/Q vssd1 vssd1 vccd1 vccd1 _11979_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13718_ _14188_/CLK _13718_/D vssd1 vssd1 vccd1 vccd1 _13718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _14139_/CLK _13649_/D vssd1 vssd1 vccd1 vccd1 _13649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07170_ _14479_/Q _07164_/X _06719_/X _07166_/X _07169_/X vssd1 vssd1 vccd1 vccd1
+ _14479_/D sky130_fd_sc_hd__o221a_1
XFILLER_199_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput602 _13259_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09811_ _13348_/Q vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__inv_2
XFILLER_173_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09742_ _10128_/A _09742_/B _09741_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__or3b_2
X_06954_ _06954_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _14574_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09673_ _14597_/Q _14594_/Q _06865_/A _06875_/Y vssd1 vssd1 vccd1 vccd1 _09673_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06885_ _06899_/A _06885_/B vssd1 vssd1 vccd1 vccd1 _14593_/D sky130_fd_sc_hd__nor2_1
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08624_ _13761_/Q _08618_/X _08534_/X _08619_/X _08620_/X vssd1 vssd1 vccd1 vccd1
+ _13761_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08555_ _13793_/Q _08552_/X _08553_/X _08554_/X _08550_/X vssd1 vssd1 vccd1 vccd1
+ _13793_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07506_ _14317_/Q _07499_/X _07330_/X _07501_/X _07503_/X vssd1 vssd1 vccd1 vccd1
+ _14317_/D sky130_fd_sc_hd__o221a_1
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08486_ _08486_/A vssd1 vssd1 vccd1 vccd1 _08486_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07437_ _14352_/Q _07432_/X _07341_/X _07433_/X _07434_/X vssd1 vssd1 vccd1 vccd1
+ _14352_/D sky130_fd_sc_hd__o221a_1
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07368_ _14381_/Q _07361_/X _07367_/X _07363_/X _07359_/X vssd1 vssd1 vccd1 vccd1
+ _14381_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09107_ _13516_/Q _09103_/X _08950_/X _09104_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _13516_/D sky130_fd_sc_hd__o221a_1
X_07299_ _14406_/Q _07238_/A _06845_/X _07240_/A _07295_/X vssd1 vssd1 vccd1 vccd1
+ _14406_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09038_ _13553_/Q _09030_/X _08954_/X _09031_/X _09036_/X vssd1 vssd1 vccd1 vccd1
+ _13553_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11000_ _13399_/Q _10804_/X _13711_/Q _10936_/X vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12951_ _12555_/X _12950_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__mux2_1
XPHY_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _13496_/Q vssd1 vssd1 vccd1 vccd1 _11902_/Y sky130_fd_sc_hd__inv_2
XPHY_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12531_/X _12881_/X _12922_/S vssd1 vssd1 vccd1 vccd1 _12882_/X sky130_fd_sc_hd__mux2_1
XANTENNA_200 _12282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 _13286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/CLK _14621_/D vssd1 vssd1 vccd1 vccd1 _14621_/Q sky130_fd_sc_hd__dfxtp_1
X_11833_ _13417_/Q _11747_/X _13736_/Q _12416_/S _11832_/X vssd1 vssd1 vccd1 vccd1
+ _11866_/B sky130_fd_sc_hd__a221oi_2
XPHY_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14552_ _14629_/CLK _14552_/D vssd1 vssd1 vccd1 vccd1 _14552_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _14358_/Q vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__inv_2
XPHY_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _14094_/CLK _13503_/D vssd1 vssd1 vccd1 vccd1 _13503_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _13510_/Q vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14483_ _14637_/CLK _14483_/D vssd1 vssd1 vccd1 vccd1 _14483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11695_/A vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13434_ _14143_/CLK _13434_/D vssd1 vssd1 vccd1 vccd1 _13434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10646_ _13431_/Q vssd1 vssd1 vccd1 vccd1 _10646_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13365_ _14639_/CLK _13365_/D vssd1 vssd1 vccd1 vccd1 _13365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10577_ _10575_/Y _10455_/X _10576_/Y _10458_/X vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12316_ _10561_/Y _14527_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13296_ _13877_/CLK _13296_/D vssd1 vssd1 vccd1 vccd1 _13296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12247_ _12247_/A vssd1 vssd1 vccd1 vccd1 _12247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ vssd1 vssd1 vccd1 vccd1 _12178_/HI _12178_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11129_ _13877_/Q vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06670_ _06667_/Y _06669_/X _06667_/Y _06669_/X vssd1 vssd1 vccd1 vccd1 _06670_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08340_ _08814_/A _08340_/B _08584_/C _08584_/D vssd1 vssd1 vccd1 vccd1 _11650_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_127_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ _08341_/A _11689_/A vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__or2_2
XFILLER_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ _07262_/A vssd1 vssd1 vccd1 vccd1 _07222_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07084_ _14521_/Q _07014_/A _07083_/X _07017_/A _07079_/X vssd1 vssd1 vccd1 vccd1
+ _14521_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput410 _12089_/LO vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput421 _12237_/A vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput432 _12247_/A vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput443 _12085_/LO vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput454 _12241_/X vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput465 _10121_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__clkbuf_2
Xoutput476 _10144_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__clkbuf_2
Xoutput487 _12119_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput498 _12129_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07986_ _08133_/A vssd1 vssd1 vccd1 vccd1 _08017_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09725_ _09717_/X _09724_/X _09717_/X _09724_/X vssd1 vssd1 vccd1 vccd1 _10140_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06937_ _06956_/A vssd1 vssd1 vccd1 vccd1 _06937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09656_ _09656_/A vssd1 vssd1 vccd1 vccd1 _09656_/Y sky130_fd_sc_hd__inv_2
X_06868_ _14596_/Q vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__inv_2
X_08607_ _13772_/Q _08599_/X _08606_/X _08601_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _13772_/D sky130_fd_sc_hd__o221a_1
XFILLER_3_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09587_ _09583_/X _09586_/X _13260_/Q _09584_/X vssd1 vssd1 vccd1 vccd1 _13228_/D
+ sky130_fd_sc_hd__o22a_1
X_06799_ _14614_/Q _06787_/X _06532_/X _08243_/A _06785_/X vssd1 vssd1 vccd1 vccd1
+ _14614_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08538_/X sky130_fd_sc_hd__clkbuf_2
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08469_ _08469_/A vssd1 vssd1 vccd1 vccd1 _08469_/X sky130_fd_sc_hd__clkbuf_2
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10500_ _11685_/A vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__buf_4
XFILLER_183_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _11478_/Y _11419_/X _11479_/Y _11421_/X vssd1 vssd1 vccd1 vccd1 _11480_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _11401_/A vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13150_ _13149_/X _12653_/X _13178_/S vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__mux2_1
X_10362_ _14485_/Q vssd1 vssd1 vccd1 vccd1 _10362_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ vssd1 vssd1 vccd1 vccd1 _12101_/HI _12101_/LO sky130_fd_sc_hd__conb_1
XFILLER_139_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10293_ _13462_/Q vssd1 vssd1 vccd1 vccd1 _10293_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13081_ _12619_/X _13080_/X _13145_/S vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12032_ _09770_/A _13146_/S _09882_/A _12954_/S vssd1 vssd1 vccd1 vccd1 _12032_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13983_ _14100_/CLK _13983_/D vssd1 vssd1 vccd1 vccd1 _13983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12934_ _12933_/X _12547_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12527_/X _12864_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14604_ _14629_/CLK _14604_/D vssd1 vssd1 vccd1 vccd1 _14604_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11816_ _13930_/Q vssd1 vssd1 vccd1 vccd1 _11816_/Y sky130_fd_sc_hd__inv_2
XPHY_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12511_/X input359/X _13080_/S vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14535_ _14538_/CLK _14535_/D vssd1 vssd1 vccd1 vccd1 _14535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11747_ _11747_/A vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__clkbuf_4
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14495_/CLK _14466_/D vssd1 vssd1 vccd1 vccd1 _14466_/Q sky130_fd_sc_hd__dfxtp_1
X_11678_ _14317_/Q vssd1 vssd1 vccd1 vccd1 _11678_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13417_ _14173_/CLK _13417_/D vssd1 vssd1 vccd1 vccd1 _13417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10629_ _10627_/Y _10484_/X _10628_/Y _10487_/X vssd1 vssd1 vccd1 vccd1 _10629_/X
+ sky130_fd_sc_hd__o22a_1
X_14397_ _14633_/CLK _14397_/D vssd1 vssd1 vccd1 vccd1 _14397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _14538_/CLK _13348_/D vssd1 vssd1 vccd1 vccd1 _13348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13279_ _14538_/CLK _13279_/D vssd1 vssd1 vccd1 vccd1 _13279_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_174_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07840_ _14154_/Q _07837_/X _07746_/X _07838_/X _07839_/X vssd1 vssd1 vccd1 vccd1
+ _14154_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07771_ _08162_/A vssd1 vssd1 vccd1 vccd1 _07771_/X sky130_fd_sc_hd__buf_4
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09510_ _12853_/S vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__clkbuf_2
X_06722_ _07712_/A vssd1 vssd1 vccd1 vccd1 _06722_/X sky130_fd_sc_hd__buf_2
XFILLER_65_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09441_ _09444_/A _12963_/X vssd1 vssd1 vccd1 vccd1 _13301_/D sky130_fd_sc_hd__and2_1
XFILLER_65_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06653_ _08981_/A _06652_/X _06632_/A _06652_/X vssd1 vssd1 vccd1 vccd1 _06653_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09372_ _09376_/A _12803_/X vssd1 vssd1 vccd1 vccd1 _13357_/D sky130_fd_sc_hd__and2_1
XFILLER_209_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06584_ input98/X vssd1 vssd1 vccd1 vccd1 _06584_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ _13908_/Q _08318_/X _08167_/X _08319_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _13908_/D sky130_fd_sc_hd__o221a_1
XFILLER_90_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ _13945_/Q _08246_/X _08171_/X _08247_/X _08249_/X vssd1 vssd1 vccd1 vccd1
+ _13945_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07205_ _07213_/A vssd1 vssd1 vccd1 vccd1 _07205_/X sky130_fd_sc_hd__buf_2
XFILLER_88_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _13979_/Q _08174_/X _08183_/X _08176_/X _08184_/X vssd1 vssd1 vccd1 vccd1
+ _13979_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07136_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07067_ _14531_/Q _07061_/X _06817_/X _07062_/X _07063_/X vssd1 vssd1 vccd1 vccd1
+ _14531_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07969_ _14085_/Q _07965_/X _07723_/X _07967_/X _07960_/X vssd1 vssd1 vccd1 vccd1
+ _14085_/D sky130_fd_sc_hd__o221a_1
XFILLER_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09708_ _14590_/Q _14586_/Q _06893_/X _06909_/Y vssd1 vssd1 vccd1 vccd1 _09708_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10976_/Y _10977_/X _10978_/Y _10979_/X vssd1 vssd1 vccd1 vccd1 _10980_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _06909_/Y _14578_/Q _14586_/Q _06938_/Y vssd1 vssd1 vccd1 vccd1 _09641_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _09821_/Y _13335_/Q _12650_/S vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__mux2_1
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _13887_/Q vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__inv_2
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12581_ _09936_/X _13306_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12581_/X sky130_fd_sc_hd__mux2_1
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14320_ _14481_/CLK _14320_/D vssd1 vssd1 vccd1 vccd1 _14320_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11532_ _14626_/Q vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__inv_2
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14251_ _14325_/CLK _14251_/D vssd1 vssd1 vccd1 vccd1 _14251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11463_ _11454_/Y _11455_/X _11456_/Y _11457_/X _11462_/X vssd1 vssd1 vccd1 vccd1
+ _11464_/D sky130_fd_sc_hd__o221a_1
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13202_ _13368_/CLK _13202_/D vssd1 vssd1 vccd1 vccd1 _13202_/Q sky130_fd_sc_hd__dfxtp_2
X_10414_ _10409_/Y _10228_/X _10410_/Y _10231_/X _10413_/X vssd1 vssd1 vccd1 vccd1
+ _10421_/C sky130_fd_sc_hd__o221a_1
XFILLER_109_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14182_ _14183_/CLK _14182_/D vssd1 vssd1 vccd1 vccd1 _14182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11394_ _11375_/X _11394_/B _11394_/C _11394_/D vssd1 vssd1 vccd1 vccd1 _11395_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _12645_/X _13132_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__mux2_1
X_10345_ _10343_/Y _10156_/X _10344_/Y _10159_/X vssd1 vssd1 vccd1 vccd1 _10345_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13064_ _12612_/X input356/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13064_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10276_ _11013_/A vssd1 vssd1 vccd1 vccd1 _10276_/X sky130_fd_sc_hd__buf_2
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _12013_/Y _10220_/A _12014_/Y _10223_/A vssd1 vssd1 vccd1 vccd1 _12015_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13966_ _14094_/CLK _13966_/D vssd1 vssd1 vccd1 vccd1 _13966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _12540_/X _12916_/X _13177_/S vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13897_ _14169_/CLK _13897_/D vssd1 vssd1 vccd1 vccd1 _13897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12848_ _12523_/X input331/X _13112_/S vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12779_ _09524_/X _12778_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13219_/D sky130_fd_sc_hd__mux2_1
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14518_ _14637_/CLK _14518_/D vssd1 vssd1 vccd1 vccd1 _14518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _14529_/CLK _14449_/D vssd1 vssd1 vccd1 vccd1 _14449_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09990_ _13366_/Q _09990_/B vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _13598_/Q _08929_/X _08940_/X _08931_/X _08938_/X vssd1 vssd1 vccd1 vccd1
+ _13598_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08872_ _13629_/Q _08868_/X _08556_/X _08869_/X _08871_/X vssd1 vssd1 vccd1 vccd1
+ _13629_/D sky130_fd_sc_hd__o221a_1
XFILLER_170_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07823_ _14164_/Q _07819_/X _07719_/X _07821_/X _07822_/X vssd1 vssd1 vccd1 vccd1
+ _14164_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07754_ _14190_/Q _07745_/X _07753_/X _07747_/X _07743_/X vssd1 vssd1 vccd1 vccd1
+ _14190_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06705_ _06695_/X _06703_/X _06704_/Y vssd1 vssd1 vccd1 vccd1 _06705_/X sky130_fd_sc_hd__o21a_1
X_07685_ _14219_/Q _07679_/X _07381_/X _07680_/X _07684_/X vssd1 vssd1 vccd1 vccd1
+ _14219_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09424_ _09426_/A _13035_/X vssd1 vssd1 vccd1 vccd1 _13315_/D sky130_fd_sc_hd__and2_1
XFILLER_168_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06636_ _08962_/A input98/X _06628_/Y _06584_/Y vssd1 vssd1 vccd1 vccd1 _06636_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09355_ _09357_/A _12879_/X vssd1 vssd1 vccd1 vccd1 _13370_/D sky130_fd_sc_hd__and2_1
XFILLER_55_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06567_ _06696_/A vssd1 vssd1 vccd1 vccd1 _06567_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ _13919_/Q _08302_/X _08140_/X _08303_/X _08305_/X vssd1 vssd1 vccd1 vccd1
+ _13919_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _09327_/A vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06498_ _06498_/A _06498_/B _06498_/C vssd1 vssd1 vccd1 vccd1 _06499_/D sky130_fd_sc_hd__or3_4
XFILLER_205_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _08246_/A vssd1 vssd1 vccd1 vccd1 _08237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ _13986_/Q _08161_/X _08167_/X _08163_/X _08159_/X vssd1 vssd1 vccd1 vccd1
+ _13986_/D sky130_fd_sc_hd__o221a_1
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07119_ _07136_/A vssd1 vssd1 vccd1 vccd1 _07119_/X sky130_fd_sc_hd__clkbuf_2
X_08099_ _08822_/A vssd1 vssd1 vccd1 vccd1 _08099_/X sky130_fd_sc_hd__buf_4
XFILLER_49_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _12440_/S sky130_fd_sc_hd__or2_1
XFILLER_66_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _10107_/A _10098_/A vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__or2_2
XFILLER_66_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13820_ _14095_/CLK _13820_/D vssd1 vssd1 vccd1 vccd1 _13820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13751_ _14110_/CLK _13751_/D vssd1 vssd1 vccd1 vccd1 _13751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10963_ _11435_/A vssd1 vssd1 vccd1 vccd1 _10963_/X sky130_fd_sc_hd__buf_2
X_12702_ _09560_/X _12701_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13682_ _14143_/CLK _13682_/D vssd1 vssd1 vccd1 vccd1 _13682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ _14106_/Q vssd1 vssd1 vccd1 vccd1 _10894_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _13328_/Q _12632_/X _12635_/S vssd1 vssd1 vccd1 vccd1 _12633_/X sky130_fd_sc_hd__mux2_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12564_ _13299_/Q _12563_/X _12651_/S vssd1 vssd1 vccd1 vccd1 _12564_/X sky130_fd_sc_hd__mux2_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _14459_/CLK _14303_/D vssd1 vssd1 vccd1 vccd1 _14303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11515_ _13410_/Q _11514_/X _13722_/Q _11408_/X vssd1 vssd1 vccd1 vccd1 _11515_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_12_1904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12495_ _12494_/X _06982_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12495_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14234_ _14611_/CLK _14234_/D vssd1 vssd1 vccd1 vccd1 _14234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11446_ _13603_/Q vssd1 vssd1 vccd1 vccd1 _11446_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14165_ _14173_/CLK _14165_/D vssd1 vssd1 vccd1 vccd1 _14165_/Q sky130_fd_sc_hd__dfxtp_1
X_11377_ _14350_/Q vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ _12637_/X input345/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10328_ _13580_/Q vssd1 vssd1 vccd1 vccd1 _10328_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14096_ _14100_/CLK _14096_/D vssd1 vssd1 vccd1 vccd1 _14096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13047_ _12602_/X _13046_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13047_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10259_ _13618_/Q vssd1 vssd1 vccd1 vccd1 _10259_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13949_ _14107_/CLK _13949_/D vssd1 vssd1 vccd1 vccd1 _13949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ _14334_/Q _07467_/X _07388_/X _07468_/X _07469_/X vssd1 vssd1 vccd1 vccd1
+ _14334_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09140_ _13499_/Q _09135_/X _08895_/X _09137_/X _09139_/X vssd1 vssd1 vccd1 vccd1
+ _13499_/D sky130_fd_sc_hd__o221a_1
X_09071_ _13537_/Q _09067_/X _08822_/X _09069_/X _09061_/X vssd1 vssd1 vccd1 vccd1
+ _13537_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08022_ _08341_/A _10201_/A vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__or2_2
XFILLER_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09973_ _09973_/A vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__inv_2
XFILLER_118_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08924_ _13604_/Q _08916_/X _08922_/X _08918_/X _08923_/X vssd1 vssd1 vccd1 vccd1
+ _13604_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08855_ _08871_/A vssd1 vssd1 vccd1 vccd1 _08855_/X sky130_fd_sc_hd__clkbuf_2
XPHY_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__inv_2
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08786_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__buf_1
XFILLER_2_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _14197_/Q _07732_/X _07736_/X _07734_/X _07730_/X vssd1 vssd1 vccd1 vccd1
+ _14197_/D sky130_fd_sc_hd__o221a_1
XPHY_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07668_ _14228_/Q _07661_/X _07358_/X _07662_/X _07666_/X vssd1 vssd1 vccd1 vccd1
+ _14228_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09407_ _09407_/A _13111_/X vssd1 vssd1 vccd1 vccd1 _13328_/D sky130_fd_sc_hd__and2_1
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06619_ input94/X _06617_/Y _06574_/Y _08979_/A vssd1 vssd1 vccd1 vccd1 _06619_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07599_ _14266_/Q _07597_/X _07362_/X _07598_/X _07593_/X vssd1 vssd1 vccd1 vccd1
+ _14266_/D sky130_fd_sc_hd__o221a_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09338_ _13384_/Q _09275_/A _08190_/A _09277_/A _09352_/A vssd1 vssd1 vccd1 vccd1
+ _13384_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _13423_/Q _09205_/A _08985_/X _09207_/A _09267_/X vssd1 vssd1 vccd1 vccd1
+ _13423_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _14309_/Q vssd1 vssd1 vccd1 vccd1 _11300_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12280_ _12072_/Y _13381_/Q _12281_/S vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _13443_/Q vssd1 vssd1 vccd1 vccd1 _11231_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162_ _13442_/Q vssd1 vssd1 vccd1 vccd1 _11162_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10113_ _10113_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _12461_/S sky130_fd_sc_hd__or2_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11093_ _13993_/Q vssd1 vssd1 vccd1 vccd1 _11093_/Y sky130_fd_sc_hd__inv_2
XPHY_7320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput310 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _06495_/A sky130_fd_sc_hd__clkbuf_1
XPHY_7331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput321 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _06497_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_1_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10044_ _13365_/Q _09988_/B _09989_/A vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__o21a_1
Xinput332 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 input332/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput343 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input343/X sky130_fd_sc_hd__buf_4
XPHY_7364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput354 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 input354/X sky130_fd_sc_hd__buf_4
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput365 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _09796_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13803_ _13996_/CLK _13803_/D vssd1 vssd1 vccd1 vccd1 _13803_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11995_ _11990_/Y _10150_/A _11991_/Y _10153_/A _11994_/X vssd1 vssd1 vccd1 vccd1
+ _12030_/A sky130_fd_sc_hd__o221a_2
XPHY_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13734_ _14169_/CLK _13734_/D vssd1 vssd1 vccd1 vccd1 _13734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _13834_/Q vssd1 vssd1 vccd1 vccd1 _10946_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _14119_/CLK _13665_/D vssd1 vssd1 vccd1 vccd1 _13665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _10875_/Y _10749_/X _10876_/Y _10751_/X vssd1 vssd1 vccd1 vccd1 _10877_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _13321_/Q _12615_/X input39/X vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13596_ _14188_/CLK _13596_/D vssd1 vssd1 vccd1 vccd1 _13596_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12547_ _13292_/Q _12546_/X _12610_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12478_ _12477_/X _06957_/Y _12505_/S vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__mux2_2
XFILLER_126_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 _10797_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14217_ _14529_/CLK _14217_/D vssd1 vssd1 vccd1 vccd1 _14217_/Q sky130_fd_sc_hd__dfxtp_1
X_11429_ _11429_/A vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__buf_2
XFILLER_12_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ _14188_/CLK _14148_/D vssd1 vssd1 vccd1 vccd1 _14148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14079_ _14305_/CLK _14079_/D vssd1 vssd1 vccd1 vccd1 _14079_/Q sky130_fd_sc_hd__dfxtp_1
X_06970_ _14569_/Q vssd1 vssd1 vccd1 vccd1 _06970_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08640_ _13752_/Q _08635_/X _08558_/X _08636_/X _08637_/X vssd1 vssd1 vccd1 vccd1
+ _13752_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08571_ _13786_/Q _08565_/X _08570_/X _08567_/X _08563_/X vssd1 vssd1 vccd1 vccd1
+ _13786_/D sky130_fd_sc_hd__o221a_1
XFILLER_110_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _14307_/Q _07516_/X _07356_/X _07517_/X _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14307_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07453_ _14344_/Q _07450_/X _07362_/X _07451_/X _07452_/X vssd1 vssd1 vccd1 vccd1
+ _14344_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07384_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09123_ _13506_/Q _09119_/X _08974_/X _09120_/X _09117_/X vssd1 vssd1 vccd1 vccd1
+ _13506_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09054_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08005_ _14063_/Q _07999_/X _07778_/X _08000_/X _08003_/X vssd1 vssd1 vccd1 vccd1
+ _14063_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09956_ _13288_/Q _13287_/Q _09883_/B vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08907_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08907_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ _09887_/A _09961_/A vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__or2_2
XFILLER_135_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08838_ _08879_/A vssd1 vssd1 vccd1 vccd1 _08871_/A sky130_fd_sc_hd__buf_2
XPHY_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _08777_/A vssd1 vssd1 vccd1 vccd1 _08769_/X sky130_fd_sc_hd__clkbuf_2
XPHY_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _13668_/Q vssd1 vssd1 vccd1 vccd1 _10800_/Y sky130_fd_sc_hd__inv_2
XPHY_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11775_/Y _11689_/X _11776_/Y _11691_/X _11779_/X vssd1 vssd1 vccd1 vccd1
+ _11781_/D sky130_fd_sc_hd__o221a_1
XPHY_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _11441_/A vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__buf_1
XPHY_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13450_ _14183_/CLK _13450_/D vssd1 vssd1 vccd1 vccd1 _13450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10662_ _10660_/Y _10462_/X _10661_/Y _10465_/X vssd1 vssd1 vccd1 vccd1 _10662_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_51_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12401_ _13220_/Q _06595_/A _12407_/S vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13381_ _14538_/CLK _13381_/D vssd1 vssd1 vccd1 vccd1 _13381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10593_ _14255_/Q vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12332_ _13195_/Q input93/X _12368_/S vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12263_ _12049_/Y _13364_/Q _12267_/S vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14002_ _14110_/CLK _14002_/D vssd1 vssd1 vccd1 vccd1 _14002_/Q sky130_fd_sc_hd__dfxtp_1
X_11214_ _14268_/Q vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12194_ vssd1 vssd1 vccd1 vccd1 _12194_/HI _12194_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11145_ _11140_/Y _10963_/X _11141_/Y _10965_/X _11144_/X vssd1 vssd1 vccd1 vccd1
+ _11158_/B sky130_fd_sc_hd__o221a_2
XFILLER_123_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _11057_/X _11076_/B _11076_/C _11076_/D vssd1 vssd1 vccd1 vccd1 _11077_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput140 la_data_in[76] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__buf_1
XPHY_7161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput151 la_data_in[86] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__buf_1
XFILLER_133_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _13381_/Q _10026_/B _10026_/Y vssd1 vssd1 vccd1 vccd1 _10027_/X sky130_fd_sc_hd__o21a_1
Xinput162 la_data_in[96] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__buf_1
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 la_oenb[105] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_hd__buf_1
XPHY_7194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 la_oenb[115] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_hd__buf_1
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 la_oenb[125] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__buf_1
XFILLER_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11978_ _14207_/Q vssd1 vssd1 vccd1 vccd1 _11978_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13717_ _14146_/CLK _13717_/D vssd1 vssd1 vccd1 vccd1 _13717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10929_ _11403_/A vssd1 vssd1 vccd1 vccd1 _10929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ _14139_/CLK _13648_/D vssd1 vssd1 vccd1 vccd1 _13648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13579_ _14173_/CLK _13579_/D vssd1 vssd1 vccd1 vccd1 _13579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput603 _13260_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09810_ _09808_/A _09808_/B _09809_/Y vssd1 vssd1 vccd1 vccd1 _09810_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09741_ _12232_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _12505_/S sky130_fd_sc_hd__nor2_8
XFILLER_98_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06953_ _06937_/X _12308_/X _06952_/Y _06939_/X vssd1 vssd1 vccd1 vccd1 _06954_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09672_ _09637_/Y _09671_/A _09637_/A _09671_/Y vssd1 vssd1 vccd1 vccd1 _09672_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06884_ _06880_/X _12289_/X _06881_/Y _06883_/X vssd1 vssd1 vccd1 vccd1 _06885_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08623_ _13762_/Q _08618_/X _08532_/X _08619_/X _08620_/X vssd1 vssd1 vccd1 vccd1
+ _13762_/D sky130_fd_sc_hd__o221a_1
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08554_ _08554_/A vssd1 vssd1 vccd1 vccd1 _08554_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07505_ _14318_/Q _07499_/X _07428_/X _07501_/X _07503_/X vssd1 vssd1 vccd1 vccd1
+ _14318_/D sky130_fd_sc_hd__o221a_1
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08485_ _08565_/A vssd1 vssd1 vccd1 vccd1 _08486_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07436_ _14353_/Q _07432_/X _07339_/X _07433_/X _07434_/X vssd1 vssd1 vccd1 vccd1
+ _14353_/D sky130_fd_sc_hd__o221a_1
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07367_ _08155_/A vssd1 vssd1 vccd1 vccd1 _07367_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09106_ _13517_/Q _09103_/X _08948_/X _09104_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _13517_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07298_ _14407_/Q _07238_/A _06843_/B _07240_/A _07295_/X vssd1 vssd1 vccd1 vccd1
+ _14407_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _13554_/Q _09030_/X _09035_/X _09031_/X _09036_/X vssd1 vssd1 vccd1 vccd1
+ _13554_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09939_ _13308_/Q _09937_/Y _09903_/B vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _12949_/X _12555_/X _12954_/S vssd1 vssd1 vccd1 vccd1 _12950_/X sky130_fd_sc_hd__mux2_1
XPHY_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11901_ _14166_/Q vssd1 vssd1 vccd1 vccd1 _11901_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12881_ _12531_/X _12880_/X _13133_/S vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__mux2_1
XPHY_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_201 _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _09451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ _14243_/Q _11830_/X _14438_/Q _11831_/X vssd1 vssd1 vccd1 vccd1 _11832_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14620_ _14621_/CLK _14620_/D vssd1 vssd1 vccd1 vccd1 _14620_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14551_ _14629_/CLK _14551_/D vssd1 vssd1 vccd1 vccd1 _14551_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _14514_/Q vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__inv_2
XPHY_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _14094_/CLK _13502_/D vssd1 vssd1 vccd1 vccd1 _13502_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _11424_/A vssd1 vssd1 vccd1 vccd1 _10714_/X sky130_fd_sc_hd__clkbuf_2
X_14482_ _14637_/CLK _14482_/D vssd1 vssd1 vccd1 vccd1 _14482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _14473_/Q vssd1 vssd1 vccd1 vccd1 _11694_/Y sky130_fd_sc_hd__inv_2
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13433_ _14143_/CLK _13433_/D vssd1 vssd1 vccd1 vccd1 _13433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _14062_/Q vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _14639_/CLK _13364_/D vssd1 vssd1 vccd1 vccd1 _13364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10576_ _14099_/Q vssd1 vssd1 vccd1 vccd1 _10576_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12315_ _10603_/Y _14528_/Q _12318_/S vssd1 vssd1 vccd1 vccd1 _12315_/X sky130_fd_sc_hd__mux2_2
XFILLER_100_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _13352_/CLK _13295_/D vssd1 vssd1 vccd1 vccd1 _13295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12246_ _12246_/A vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12177_ vssd1 vssd1 vccd1 vccd1 _12177_/HI _12177_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ _13760_/Q vssd1 vssd1 vccd1 vccd1 _11128_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ _14343_/Q vssd1 vssd1 vccd1 vccd1 _11059_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08270_ _08411_/A _08890_/B _08744_/C _08584_/D vssd1 vssd1 vccd1 vccd1 _11689_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_127_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07221_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07262_/A sky130_fd_sc_hd__buf_2
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07152_ _14485_/Q _07092_/A _06843_/B _07094_/A _07147_/X vssd1 vssd1 vccd1 vccd1
+ _14485_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07083_ _08268_/A vssd1 vssd1 vccd1 vccd1 _07083_/X sky130_fd_sc_hd__buf_2
Xoutput400 _12200_/X vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__clkbuf_2
Xoutput411 _12090_/LO vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput422 _12238_/A vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput433 _12248_/A vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput444 _12096_/LO vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput455 _12242_/X vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__clkbuf_2
Xoutput466 _10123_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput477 _10146_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__clkbuf_2
Xoutput488 _12120_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput499 _12130_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _14075_/Q _07982_/X _07749_/X _07983_/X _07978_/X vssd1 vssd1 vccd1 vccd1
+ _14075_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09724_ _09720_/X _09723_/X _09720_/X _09723_/X vssd1 vssd1 vccd1 vccd1 _09724_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06936_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06954_/A sky130_fd_sc_hd__buf_2
XFILLER_5_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09655_ _06893_/A _14582_/Q _14590_/Q _06924_/Y vssd1 vssd1 vccd1 vccd1 _09656_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_3_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06867_ _06877_/A _06867_/B vssd1 vssd1 vccd1 vccd1 _14597_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08606_ _09009_/A vssd1 vssd1 vccd1 vccd1 _08606_/X sky130_fd_sc_hd__buf_4
X_09586_ _09586_/A _12331_/X vssd1 vssd1 vccd1 vccd1 _09586_/X sky130_fd_sc_hd__and2_2
XFILLER_93_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06798_ _09035_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__buf_4
X_08537_ _08645_/A vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__clkbuf_4
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _08468_/A vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__clkbuf_2
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07419_ _14361_/Q _07411_/X _07315_/X _07414_/X _07415_/X vssd1 vssd1 vccd1 vccd1
+ _14361_/D sky130_fd_sc_hd__o221a_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08399_ _13865_/Q _08396_/X _08259_/X _08397_/X _08392_/X vssd1 vssd1 vccd1 vccd1
+ _13865_/D sky130_fd_sc_hd__o221a_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10430_ _11637_/A vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10361_ _13194_/Q _10276_/X _14017_/Q _10203_/X _10360_/X vssd1 vssd1 vccd1 vccd1
+ _10361_/X sky130_fd_sc_hd__a221o_2
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12100_ vssd1 vssd1 vccd1 vccd1 _12100_/HI _12100_/LO sky130_fd_sc_hd__conb_1
XFILLER_191_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13080_ _12619_/X input330/X _13080_/S vssd1 vssd1 vccd1 vccd1 _13080_/X sky130_fd_sc_hd__mux2_1
X_10292_ _14132_/Q vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ _09770_/B _13146_/S _09882_/B _12954_/S vssd1 vssd1 vccd1 vccd1 _12031_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_137_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13982_ _14100_/CLK _13982_/D vssd1 vssd1 vccd1 vccd1 _13982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12933_ _12547_/X _12932_/X _13113_/S vssd1 vssd1 vccd1 vccd1 _12933_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12527_/X input344/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14633_/CLK _14603_/D vssd1 vssd1 vccd1 vccd1 _14603_/Q sky130_fd_sc_hd__dfxtp_1
X_11815_ _11810_/Y _11679_/X _11811_/Y _11681_/X _11814_/X vssd1 vssd1 vccd1 vccd1
+ _11822_/C sky130_fd_sc_hd__o221a_1
XPHY_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _09537_/X _12794_/X _13179_/S vssd1 vssd1 vccd1 vccd1 _13215_/D sky130_fd_sc_hd__mux2_1
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _11741_/Y _11633_/X _11742_/Y _11635_/X _11745_/X vssd1 vssd1 vccd1 vccd1
+ _11782_/A sky130_fd_sc_hd__o221a_1
X_14534_ _14611_/CLK _14534_/D vssd1 vssd1 vccd1 vccd1 _14534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11677_ _11668_/Y _11669_/X _11670_/Y _11671_/X _11676_/X vssd1 vssd1 vccd1 vccd1
+ _11698_/B sky130_fd_sc_hd__o221a_2
X_14465_ _14595_/CLK _14465_/D vssd1 vssd1 vccd1 vccd1 _14465_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13416_ _14178_/CLK _13416_/D vssd1 vssd1 vccd1 vccd1 _13416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10628_ _14373_/Q vssd1 vssd1 vccd1 vccd1 _10628_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14396_ _14629_/CLK _14396_/D vssd1 vssd1 vccd1 vccd1 _14396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13347_ _14538_/CLK _13347_/D vssd1 vssd1 vccd1 vccd1 _13347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10559_ _10554_/Y _10506_/X _10555_/Y _10509_/X _10558_/X vssd1 vssd1 vccd1 vccd1
+ _10560_/D sky130_fd_sc_hd__o221a_1
Xclkbuf_2_1_0_register_file.clk_i clkbuf_0_register_file.clk_i/X vssd1 vssd1 vccd1
+ vccd1 _13370_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13278_ _14573_/CLK _13278_/D vssd1 vssd1 vccd1 vccd1 _13278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_170_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12229_ _12231_/A vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07770_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06721_ _08827_/A vssd1 vssd1 vccd1 vccd1 _07712_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09440_ _09444_/A _12959_/X vssd1 vssd1 vccd1 vccd1 _13302_/D sky130_fd_sc_hd__and2_1
X_06652_ _06542_/X _09051_/A _06542_/X _09051_/A vssd1 vssd1 vccd1 vccd1 _06652_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09371_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06583_ input98/X vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08322_ _13909_/Q _08318_/X _08165_/X _08319_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _13909_/D sky130_fd_sc_hd__o221a_1
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08253_ _13946_/Q _08246_/X _08169_/X _08247_/X _08249_/X vssd1 vssd1 vccd1 vccd1
+ _13946_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07204_ _14460_/Q _07201_/X _06793_/X _07202_/X _07197_/X vssd1 vssd1 vccd1 vccd1
+ _14460_/D sky130_fd_sc_hd__o221a_1
X_08184_ _08184_/A vssd1 vssd1 vccd1 vccd1 _08184_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07135_ _14496_/Q _07127_/X _06801_/X _07128_/X _07131_/X vssd1 vssd1 vccd1 vccd1
+ _14496_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07066_ _14532_/Q _07061_/X _06814_/X _07062_/X _07063_/X vssd1 vssd1 vccd1 vccd1
+ _14532_/D sky130_fd_sc_hd__o221a_1
XFILLER_121_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _14086_/Q _07965_/X _07719_/X _07967_/X _07960_/X vssd1 vssd1 vccd1 vccd1
+ _14086_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09707_ _14570_/Q _14569_/Q _06967_/Y _06970_/Y vssd1 vssd1 vccd1 vccd1 _09707_/X
+ sky130_fd_sc_hd__o22a_1
X_06919_ _06956_/A vssd1 vssd1 vccd1 vccd1 _06919_/X sky130_fd_sc_hd__buf_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ _14123_/Q _07892_/X _07825_/X _07894_/X _07897_/X vssd1 vssd1 vccd1 vccd1
+ _14123_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _14588_/Q _14580_/Q _06902_/Y _06930_/Y vssd1 vssd1 vccd1 vccd1 _09640_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _09573_/A _12361_/X vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__and2_1
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _13770_/Q vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__inv_2
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12580_ _13307_/Q _12579_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__mux2_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11531_ _14353_/Q vssd1 vssd1 vccd1 vccd1 _11531_/Y sky130_fd_sc_hd__inv_2
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14250_ _14325_/CLK _14250_/D vssd1 vssd1 vccd1 vccd1 _14250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11462_ _11458_/Y _11459_/X _11460_/Y _11461_/X vssd1 vssd1 vccd1 vccd1 _11462_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13368_/CLK _13201_/D vssd1 vssd1 vccd1 vccd1 _13201_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _10411_/Y _10234_/X _10412_/Y _10237_/X vssd1 vssd1 vccd1 vccd1 _10413_/X
+ sky130_fd_sc_hd__o22a_1
X_14181_ _14183_/CLK _14181_/D vssd1 vssd1 vccd1 vccd1 _14181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11393_ _11388_/Y _11219_/X _11389_/Y _11221_/X _11392_/X vssd1 vssd1 vccd1 vccd1
+ _11394_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13132_ _12645_/X input340/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_1
X_10344_ _13620_/Q vssd1 vssd1 vccd1 vccd1 _10344_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ _12610_/X _13062_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13063_/X sky130_fd_sc_hd__mux2_1
X_10275_ _11485_/A vssd1 vssd1 vccd1 vccd1 _11013_/A sky130_fd_sc_hd__buf_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _14403_/Q vssd1 vssd1 vccd1 vccd1 _12014_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13965_ _14094_/CLK _13965_/D vssd1 vssd1 vccd1 vccd1 _13965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12916_ _12540_/X input347/X _13176_/S vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13896_ _14130_/CLK _13896_/D vssd1 vssd1 vccd1 vccd1 _13896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12847_ _12522_/X _12846_/X _13099_/S vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12778_ _09524_/X _12777_/X _12794_/S vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14517_ _14637_/CLK _14517_/D vssd1 vssd1 vccd1 vccd1 _14517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11729_ _14201_/Q vssd1 vssd1 vccd1 vccd1 _11729_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14448_ _14529_/CLK _14448_/D vssd1 vssd1 vccd1 vccd1 _14448_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14379_ _14627_/CLK _14379_/D vssd1 vssd1 vccd1 vccd1 _14379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08940_ _08940_/A vssd1 vssd1 vccd1 vccd1 _08940_/X sky130_fd_sc_hd__buf_6
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08871_ _08871_/A vssd1 vssd1 vccd1 vccd1 _08871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater700 _13145_/S vssd1 vssd1 vccd1 vccd1 _13141_/S sky130_fd_sc_hd__buf_8
XFILLER_6_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07822_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07753_ _08144_/A vssd1 vssd1 vccd1 vccd1 _07753_/X sky130_fd_sc_hd__buf_6
XFILLER_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06704_ _06853_/A _09035_/A _06695_/X vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__o21ai_1
X_07684_ _07715_/A vssd1 vssd1 vccd1 vccd1 _07684_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09423_ _09426_/A _13031_/X vssd1 vssd1 vccd1 vccd1 _13316_/D sky130_fd_sc_hd__and2_1
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06635_ input99/X vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__buf_2
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _09357_/A _12875_/X vssd1 vssd1 vccd1 vccd1 _13371_/D sky130_fd_sc_hd__and2_1
XFILLER_94_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06566_ _06535_/A _06564_/Y _06535_/Y _08925_/A vssd1 vssd1 vccd1 vccd1 _06566_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08305_ _08329_/A vssd1 vssd1 vccd1 vccd1 _08305_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09285_ _09318_/A vssd1 vssd1 vccd1 vccd1 _09285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06497_ _06497_/A _06497_/B _06497_/C input317/X vssd1 vssd1 vccd1 vccd1 _06498_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _13955_/Q _08229_/X _08146_/X _08230_/X _08231_/X vssd1 vssd1 vccd1 vccd1
+ _13955_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08167_ _08167_/A vssd1 vssd1 vccd1 vccd1 _08167_/X sky130_fd_sc_hd__buf_4
XFILLER_68_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07118_ _14506_/Q _07111_/X _06766_/X _07112_/X _07114_/X vssd1 vssd1 vccd1 vccd1
+ _14506_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08098_ _14013_/Q _08095_/X _07809_/X _08097_/X _08089_/X vssd1 vssd1 vccd1 vccd1
+ _14013_/D sky130_fd_sc_hd__o221a_1
XFILLER_84_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07049_ _14542_/Q _07044_/X _06778_/X _07045_/X _07046_/X vssd1 vssd1 vccd1 vccd1
+ _14542_/D sky130_fd_sc_hd__o221a_1
XFILLER_157_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10060_ _10060_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__or2_1
XPHY_7513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_6889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13750_ _14110_/CLK _13750_/D vssd1 vssd1 vccd1 vccd1 _13750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _14497_/Q vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12701_ _09560_/X _12700_/X _13141_/S vssd1 vssd1 vccd1 vccd1 _12701_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13681_ _14143_/CLK _13681_/D vssd1 vssd1 vccd1 vccd1 _13681_/Q sky130_fd_sc_hd__dfxtp_1
X_10893_ _13833_/Q vssd1 vssd1 vccd1 vccd1 _10893_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _09836_/X _13328_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12632_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12563_ _09950_/Y _13299_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12563_/X sky130_fd_sc_hd__mux2_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _11514_/A vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14302_ _14459_/CLK _14302_/D vssd1 vssd1 vccd1 vccd1 _14302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12494_ _12509_/X _06982_/Y _12494_/S vssd1 vssd1 vccd1 vccd1 _12494_/X sky130_fd_sc_hd__mux2_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_1792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11445_ _11445_/A vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__clkbuf_2
X_14233_ _14611_/CLK _14233_/D vssd1 vssd1 vccd1 vccd1 _14233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14164_ _14291_/CLK _14164_/D vssd1 vssd1 vccd1 vccd1 _14164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11376_ _14506_/Q vssd1 vssd1 vccd1 vccd1 _11376_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10327_ _14289_/Q vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13115_ _12635_/X _13114_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__mux2_1
X_14095_ _14095_/CLK _14095_/D vssd1 vssd1 vccd1 vccd1 _14095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13046_ _13045_/X _12602_/X _13050_/S vssd1 vssd1 vccd1 vccd1 _13046_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _13657_/Q vssd1 vssd1 vccd1 vccd1 _10258_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10189_ _14092_/Q vssd1 vssd1 vccd1 vccd1 _10189_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13948_ _14107_/CLK _13948_/D vssd1 vssd1 vccd1 vccd1 _13948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13879_ _13996_/CLK _13879_/D vssd1 vssd1 vccd1 vccd1 _13879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09070_ _13538_/Q _09067_/X _08895_/X _09069_/X _09061_/X vssd1 vssd1 vccd1 vccd1
+ _13538_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _09131_/A _09063_/B _09063_/C _08673_/D vssd1 vssd1 vccd1 vccd1 _10201_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_159_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09972_ _13357_/Q _09972_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08923_ _08923_/A vssd1 vssd1 vccd1 vccd1 _08923_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08854_ _13640_/Q _08852_/X _08527_/X _08853_/X _08847_/X vssd1 vssd1 vccd1 vccd1
+ _13640_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _07952_/A _11691_/A vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__or2_2
XFILLER_79_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _08879_/A vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__clkbuf_4
XPHY_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _08126_/A vssd1 vssd1 vccd1 vccd1 _07736_/X sky130_fd_sc_hd__buf_4
XPHY_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07667_ _14229_/Q _07661_/X _07356_/X _07662_/X _07666_/X vssd1 vssd1 vccd1 vccd1
+ _14229_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _09407_/A _13107_/X vssd1 vssd1 vccd1 vccd1 _13329_/D sky130_fd_sc_hd__and2_1
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06618_ input93/X vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_201_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07598_ _07606_/A vssd1 vssd1 vccd1 vccd1 _07598_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _09509_/A vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__buf_6
X_06549_ _06537_/X _06548_/X _06537_/X _06548_/X vssd1 vssd1 vccd1 vccd1 _06740_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09268_ _13424_/Q _09205_/A _08983_/X _09207_/A _09267_/X vssd1 vssd1 vccd1 vccd1
+ _13424_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08219_ _13966_/Q _08211_/X _08117_/X _08213_/X _08214_/X vssd1 vssd1 vccd1 vccd1
+ _13966_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ _13462_/Q _09135_/A _08985_/X _09137_/A _09196_/X vssd1 vssd1 vccd1 vccd1
+ _13462_/D sky130_fd_sc_hd__o221a_1
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _14074_/Q vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11161_ _11397_/A vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__buf_2
XFILLER_1_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__or2_1
XFILLER_175_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11092_ _11090_/Y _10947_/X _11091_/Y _10949_/X vssd1 vssd1 vccd1 vccd1 _11092_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_7310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput300 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _06502_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput311 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _06495_/D sky130_fd_sc_hd__clkbuf_1
XPHY_7332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ _13364_/Q _09986_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput322 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _06500_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput333 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 input333/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput344 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 input344/X sky130_fd_sc_hd__buf_6
XPHY_7365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput355 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input355/X sky130_fd_sc_hd__buf_4
XPHY_7376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput366 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _06488_/A sky130_fd_sc_hd__clkbuf_2
XPHY_7387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13802_ _13996_/CLK _13802_/D vssd1 vssd1 vccd1 vccd1 _13802_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _11992_/Y _10156_/A _11993_/Y _10159_/A vssd1 vssd1 vccd1 vccd1 _11994_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13733_ _14056_/CLK _13733_/D vssd1 vssd1 vccd1 vccd1 _13733_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10945_ _10941_/Y _10942_/X _10943_/Y _10944_/X vssd1 vssd1 vccd1 vccd1 _10945_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13664_ _14047_/CLK _13664_/D vssd1 vssd1 vccd1 vccd1 _13664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876_ _14456_/Q vssd1 vssd1 vccd1 vccd1 _10876_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _09849_/Y _13321_/Q _12634_/S vssd1 vssd1 vccd1 vccd1 _12615_/X sky130_fd_sc_hd__mux2_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _14188_/CLK _13595_/D vssd1 vssd1 vccd1 vccd1 _13595_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12546_ _09962_/Y _13292_/Q _12601_/S vssd1 vssd1 vccd1 vccd1 _12546_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12477_ _12476_/X _06957_/Y _12603_/S vssd1 vssd1 vccd1 vccd1 _12477_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_4 _10921_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14529_/CLK _14216_/D vssd1 vssd1 vccd1 vccd1 _14216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11428_ _11411_/Y _11412_/X _11417_/X _11422_/X _11427_/X vssd1 vssd1 vccd1 vccd1
+ _11465_/C sky130_fd_sc_hd__o2111a_4
XFILLER_103_1896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11359_ _11357_/Y _11165_/X _11358_/Y _11167_/X vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14147_ _14188_/CLK _14147_/D vssd1 vssd1 vccd1 vccd1 _14147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14078_ _14305_/CLK _14078_/D vssd1 vssd1 vccd1 vccd1 _14078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13029_ _12594_/X _13028_/X _13121_/S vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08570_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08570_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_208_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07521_ _14308_/Q _07516_/X _07354_/X _07517_/X _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14308_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07452_ _07476_/A vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07383_ _08171_/A vssd1 vssd1 vccd1 vccd1 _07383_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _13507_/Q _09119_/X _09051_/X _09120_/X _09117_/X vssd1 vssd1 vccd1 vccd1
+ _13507_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _13545_/Q _09048_/X _08974_/X _09049_/X _09045_/X vssd1 vssd1 vccd1 vccd1
+ _13545_/D sky130_fd_sc_hd__o221a_1
XFILLER_191_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08004_ _14064_/Q _07999_/X _07776_/X _08000_/X _08003_/X vssd1 vssd1 vccd1 vccd1
+ _14064_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09955_ _13287_/Q _12601_/S _09882_/B _12232_/A vssd1 vssd1 vccd1 vccd1 _09955_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _08971_/A vssd1 vssd1 vccd1 vccd1 _08958_/A sky130_fd_sc_hd__buf_4
XFILLER_24_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09886_ _09886_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__or2_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08837_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08837_/X sky130_fd_sc_hd__buf_4
XPHY_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08793_/A vssd1 vssd1 vccd1 vccd1 _08768_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07719_ _07719_/A vssd1 vssd1 vccd1 vccd1 _07719_/X sky130_fd_sc_hd__buf_4
XPHY_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08699_ _08723_/A vssd1 vssd1 vccd1 vccd1 _08699_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _14375_/Q vssd1 vssd1 vccd1 vccd1 _10730_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _13509_/Q vssd1 vssd1 vccd1 vccd1 _10661_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _12399_/X _13221_/Q _12655_/S vssd1 vssd1 vccd1 vccd1 _12400_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ _14538_/CLK _13380_/D vssd1 vssd1 vccd1 vccd1 _13380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10592_ _14177_/Q vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12331_ _12330_/X _13196_/Q _12647_/S vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12262_ _12048_/Y _13363_/Q _12262_/S vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _14110_/CLK _14001_/D vssd1 vssd1 vccd1 vccd1 _14001_/Q sky130_fd_sc_hd__dfxtp_1
X_11213_ _11449_/A vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__clkbuf_2
X_12193_ vssd1 vssd1 vccd1 vccd1 _12193_/HI _12193_/LO sky130_fd_sc_hd__conb_1
X_11144_ _11142_/Y _10967_/X _11143_/Y _10969_/X vssd1 vssd1 vccd1 vccd1 _11144_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11075_ _11070_/Y _10983_/X _11071_/Y _10985_/X _11074_/X vssd1 vssd1 vccd1 vccd1
+ _11076_/D sky130_fd_sc_hd__o221a_1
XPHY_7140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput130 la_data_in[67] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__buf_1
XPHY_7151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput141 la_data_in[77] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10026_ _13381_/Q _10026_/B vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__nand2_1
Xinput152 la_data_in[87] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_1
XPHY_7173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput163 la_data_in[97] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__buf_1
XFILLER_37_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput174 la_oenb[106] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_hd__buf_1
XPHY_7195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput185 la_oenb[116] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_1
XPHY_6461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput196 la_oenb[126] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__buf_1
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _13615_/Q vssd1 vssd1 vccd1 vccd1 _11977_/Y sky130_fd_sc_hd__inv_2
XPHY_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13716_ _14188_/CLK _13716_/D vssd1 vssd1 vccd1 vccd1 _13716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10928_ _13632_/Q vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13647_ _14139_/CLK _13647_/D vssd1 vssd1 vccd1 vccd1 _13647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10859_ _13552_/Q _10720_/X _13793_/Q _10721_/X vssd1 vssd1 vccd1 vccd1 _10859_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13578_ _14173_/CLK _13578_/D vssd1 vssd1 vccd1 vccd1 _13578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12529_ _13371_/Q _10034_/X _12645_/S vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput604 _13261_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09740_ _10107_/A _10090_/A vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__or2_4
X_06952_ _14574_/Q vssd1 vssd1 vccd1 vccd1 _06952_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
.ends

