magic
tech sky130A
timestamp 1638948812
<< nmos >>
rect 53 142 71 242
<< ndiff >>
rect 3 229 53 242
rect 3 211 20 229
rect 37 211 53 229
rect 3 173 53 211
rect 3 155 20 173
rect 37 155 53 173
rect 3 142 53 155
rect 71 229 121 242
rect 71 211 87 229
rect 104 211 121 229
rect 71 173 121 211
rect 71 155 87 173
rect 104 155 121 173
rect 71 142 121 155
<< ndiffc >>
rect 20 211 37 229
rect 20 155 37 173
rect 87 211 104 229
rect 87 155 104 173
<< poly >>
rect 45 282 79 290
rect 45 264 53 282
rect 71 264 79 282
rect 45 256 79 264
rect 53 242 71 256
rect 53 128 71 142
rect 45 120 79 128
rect 45 102 53 120
rect 71 102 79 120
rect 45 94 79 102
<< polycont >>
rect 53 264 71 282
rect 53 102 71 120
<< locali >>
rect 45 282 79 290
rect 45 264 53 282
rect 71 264 79 282
rect 45 256 79 264
rect 10 229 46 238
rect 10 211 20 229
rect 37 211 46 229
rect 10 202 46 211
rect 78 229 114 238
rect 78 211 87 229
rect 104 211 114 229
rect 78 202 114 211
rect 10 173 46 182
rect 10 155 20 173
rect 37 155 46 173
rect 10 146 46 155
rect 78 173 114 182
rect 78 155 87 173
rect 104 155 114 173
rect 78 146 114 155
rect 45 120 79 128
rect 45 102 53 120
rect 71 102 79 120
rect 45 94 79 102
<< labels >>
rlabel locali 62 94 62 94 1 Gate
port 1 n
rlabel locali 61 289 61 289 5 Gate
port 2 s
rlabel locali 12 162 12 162 1 Drain
port 4 n
rlabel locali 111 219 111 219 1 Source
port 5 n
rlabel locali 110 162 110 162 1 Source
port 6 n
rlabel locali 14 219 14 219 1 Drain
port 3 n
<< end >>
