VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openram_testchip
  CLASS BLOCK ;
  FOREIGN openram_testchip ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 800.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 796.000 280.970 800.000 ;
    END
  END clock
  PIN io_gpio_packet[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END io_gpio_packet[0]
  PIN io_gpio_packet[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END io_gpio_packet[10]
  PIN io_gpio_packet[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_gpio_packet[11]
  PIN io_gpio_packet[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END io_gpio_packet[12]
  PIN io_gpio_packet[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END io_gpio_packet[13]
  PIN io_gpio_packet[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 796.000 177.470 800.000 ;
    END
  END io_gpio_packet[14]
  PIN io_gpio_packet[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_gpio_packet[15]
  PIN io_gpio_packet[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_gpio_packet[16]
  PIN io_gpio_packet[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END io_gpio_packet[17]
  PIN io_gpio_packet[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 714.040 500.000 714.640 ;
    END
  END io_gpio_packet[18]
  PIN io_gpio_packet[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END io_gpio_packet[19]
  PIN io_gpio_packet[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END io_gpio_packet[1]
  PIN io_gpio_packet[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END io_gpio_packet[20]
  PIN io_gpio_packet[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.840 500.000 160.440 ;
    END
  END io_gpio_packet[21]
  PIN io_gpio_packet[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 676.640 500.000 677.240 ;
    END
  END io_gpio_packet[22]
  PIN io_gpio_packet[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_gpio_packet[23]
  PIN io_gpio_packet[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 615.440 500.000 616.040 ;
    END
  END io_gpio_packet[24]
  PIN io_gpio_packet[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END io_gpio_packet[25]
  PIN io_gpio_packet[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END io_gpio_packet[26]
  PIN io_gpio_packet[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END io_gpio_packet[27]
  PIN io_gpio_packet[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 796.000 85.470 800.000 ;
    END
  END io_gpio_packet[28]
  PIN io_gpio_packet[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END io_gpio_packet[29]
  PIN io_gpio_packet[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END io_gpio_packet[2]
  PIN io_gpio_packet[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 796.000 257.970 800.000 ;
    END
  END io_gpio_packet[30]
  PIN io_gpio_packet[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END io_gpio_packet[31]
  PIN io_gpio_packet[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_gpio_packet[32]
  PIN io_gpio_packet[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io_gpio_packet[33]
  PIN io_gpio_packet[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_gpio_packet[34]
  PIN io_gpio_packet[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END io_gpio_packet[35]
  PIN io_gpio_packet[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 796.000 55.570 800.000 ;
    END
  END io_gpio_packet[36]
  PIN io_gpio_packet[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END io_gpio_packet[37]
  PIN io_gpio_packet[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 796.000 39.470 800.000 ;
    END
  END io_gpio_packet[38]
  PIN io_gpio_packet[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 796.000 432.770 800.000 ;
    END
  END io_gpio_packet[39]
  PIN io_gpio_packet[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 796.000 352.270 800.000 ;
    END
  END io_gpio_packet[3]
  PIN io_gpio_packet[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END io_gpio_packet[40]
  PIN io_gpio_packet[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_gpio_packet[41]
  PIN io_gpio_packet[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.840 500.000 245.440 ;
    END
  END io_gpio_packet[42]
  PIN io_gpio_packet[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 513.440 500.000 514.040 ;
    END
  END io_gpio_packet[43]
  PIN io_gpio_packet[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END io_gpio_packet[44]
  PIN io_gpio_packet[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END io_gpio_packet[45]
  PIN io_gpio_packet[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END io_gpio_packet[46]
  PIN io_gpio_packet[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 727.640 500.000 728.240 ;
    END
  END io_gpio_packet[47]
  PIN io_gpio_packet[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_gpio_packet[48]
  PIN io_gpio_packet[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 796.000 446.570 800.000 ;
    END
  END io_gpio_packet[49]
  PIN io_gpio_packet[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 796.000 147.570 800.000 ;
    END
  END io_gpio_packet[4]
  PIN io_gpio_packet[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END io_gpio_packet[50]
  PIN io_gpio_packet[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_gpio_packet[51]
  PIN io_gpio_packet[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 796.000 389.070 800.000 ;
    END
  END io_gpio_packet[52]
  PIN io_gpio_packet[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 796.000 391.370 800.000 ;
    END
  END io_gpio_packet[53]
  PIN io_gpio_packet[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END io_gpio_packet[54]
  PIN io_gpio_packet[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 557.640 500.000 558.240 ;
    END
  END io_gpio_packet[55]
  PIN io_gpio_packet[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 3.440 500.000 4.040 ;
    END
  END io_gpio_packet[5]
  PIN io_gpio_packet[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END io_gpio_packet[6]
  PIN io_gpio_packet[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 796.000 306.270 800.000 ;
    END
  END io_gpio_packet[7]
  PIN io_gpio_packet[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END io_gpio_packet[8]
  PIN io_gpio_packet[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END io_gpio_packet[9]
  PIN io_in_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END io_in_select
  PIN io_logical_analyzer_packet[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 796.000 490.270 800.000 ;
    END
  END io_logical_analyzer_packet[0]
  PIN io_logical_analyzer_packet[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END io_logical_analyzer_packet[10]
  PIN io_logical_analyzer_packet[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_logical_analyzer_packet[11]
  PIN io_logical_analyzer_packet[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END io_logical_analyzer_packet[12]
  PIN io_logical_analyzer_packet[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END io_logical_analyzer_packet[13]
  PIN io_logical_analyzer_packet[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 796.000 216.570 800.000 ;
    END
  END io_logical_analyzer_packet[14]
  PIN io_logical_analyzer_packet[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END io_logical_analyzer_packet[15]
  PIN io_logical_analyzer_packet[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END io_logical_analyzer_packet[16]
  PIN io_logical_analyzer_packet[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END io_logical_analyzer_packet[17]
  PIN io_logical_analyzer_packet[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END io_logical_analyzer_packet[18]
  PIN io_logical_analyzer_packet[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END io_logical_analyzer_packet[19]
  PIN io_logical_analyzer_packet[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END io_logical_analyzer_packet[1]
  PIN io_logical_analyzer_packet[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_logical_analyzer_packet[20]
  PIN io_logical_analyzer_packet[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 796.000 425.870 800.000 ;
    END
  END io_logical_analyzer_packet[21]
  PIN io_logical_analyzer_packet[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END io_logical_analyzer_packet[22]
  PIN io_logical_analyzer_packet[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 527.040 500.000 527.640 ;
    END
  END io_logical_analyzer_packet[23]
  PIN io_logical_analyzer_packet[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END io_logical_analyzer_packet[24]
  PIN io_logical_analyzer_packet[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_logical_analyzer_packet[25]
  PIN io_logical_analyzer_packet[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_logical_analyzer_packet[26]
  PIN io_logical_analyzer_packet[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 139.440 500.000 140.040 ;
    END
  END io_logical_analyzer_packet[27]
  PIN io_logical_analyzer_packet[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END io_logical_analyzer_packet[28]
  PIN io_logical_analyzer_packet[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END io_logical_analyzer_packet[29]
  PIN io_logical_analyzer_packet[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 796.000 308.570 800.000 ;
    END
  END io_logical_analyzer_packet[2]
  PIN io_logical_analyzer_packet[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END io_logical_analyzer_packet[30]
  PIN io_logical_analyzer_packet[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_logical_analyzer_packet[31]
  PIN io_logical_analyzer_packet[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_logical_analyzer_packet[32]
  PIN io_logical_analyzer_packet[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_logical_analyzer_packet[33]
  PIN io_logical_analyzer_packet[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 796.000 101.570 800.000 ;
    END
  END io_logical_analyzer_packet[34]
  PIN io_logical_analyzer_packet[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 796.000 481.070 800.000 ;
    END
  END io_logical_analyzer_packet[35]
  PIN io_logical_analyzer_packet[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 796.000 366.070 800.000 ;
    END
  END io_logical_analyzer_packet[36]
  PIN io_logical_analyzer_packet[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 796.000 16.470 800.000 ;
    END
  END io_logical_analyzer_packet[37]
  PIN io_logical_analyzer_packet[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END io_logical_analyzer_packet[38]
  PIN io_logical_analyzer_packet[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 796.000 191.270 800.000 ;
    END
  END io_logical_analyzer_packet[39]
  PIN io_logical_analyzer_packet[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END io_logical_analyzer_packet[3]
  PIN io_logical_analyzer_packet[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_logical_analyzer_packet[40]
  PIN io_logical_analyzer_packet[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 30.640 500.000 31.240 ;
    END
  END io_logical_analyzer_packet[41]
  PIN io_logical_analyzer_packet[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 796.000 407.470 800.000 ;
    END
  END io_logical_analyzer_packet[42]
  PIN io_logical_analyzer_packet[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END io_logical_analyzer_packet[43]
  PIN io_logical_analyzer_packet[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END io_logical_analyzer_packet[44]
  PIN io_logical_analyzer_packet[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 796.000 331.570 800.000 ;
    END
  END io_logical_analyzer_packet[45]
  PIN io_logical_analyzer_packet[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END io_logical_analyzer_packet[46]
  PIN io_logical_analyzer_packet[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 796.000 27.970 800.000 ;
    END
  END io_logical_analyzer_packet[47]
  PIN io_logical_analyzer_packet[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END io_logical_analyzer_packet[48]
  PIN io_logical_analyzer_packet[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END io_logical_analyzer_packet[49]
  PIN io_logical_analyzer_packet[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 796.000 370.670 800.000 ;
    END
  END io_logical_analyzer_packet[4]
  PIN io_logical_analyzer_packet[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END io_logical_analyzer_packet[50]
  PIN io_logical_analyzer_packet[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END io_logical_analyzer_packet[51]
  PIN io_logical_analyzer_packet[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 796.000 485.670 800.000 ;
    END
  END io_logical_analyzer_packet[52]
  PIN io_logical_analyzer_packet[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END io_logical_analyzer_packet[53]
  PIN io_logical_analyzer_packet[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END io_logical_analyzer_packet[54]
  PIN io_logical_analyzer_packet[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_logical_analyzer_packet[55]
  PIN io_logical_analyzer_packet[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 796.000 138.370 800.000 ;
    END
  END io_logical_analyzer_packet[56]
  PIN io_logical_analyzer_packet[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END io_logical_analyzer_packet[57]
  PIN io_logical_analyzer_packet[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 523.640 500.000 524.240 ;
    END
  END io_logical_analyzer_packet[58]
  PIN io_logical_analyzer_packet[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 418.240 500.000 418.840 ;
    END
  END io_logical_analyzer_packet[59]
  PIN io_logical_analyzer_packet[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 796.000 294.770 800.000 ;
    END
  END io_logical_analyzer_packet[5]
  PIN io_logical_analyzer_packet[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 34.040 500.000 34.640 ;
    END
  END io_logical_analyzer_packet[60]
  PIN io_logical_analyzer_packet[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END io_logical_analyzer_packet[61]
  PIN io_logical_analyzer_packet[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 796.000 225.770 800.000 ;
    END
  END io_logical_analyzer_packet[62]
  PIN io_logical_analyzer_packet[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 666.440 500.000 667.040 ;
    END
  END io_logical_analyzer_packet[63]
  PIN io_logical_analyzer_packet[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END io_logical_analyzer_packet[64]
  PIN io_logical_analyzer_packet[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_logical_analyzer_packet[65]
  PIN io_logical_analyzer_packet[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 796.000 73.970 800.000 ;
    END
  END io_logical_analyzer_packet[66]
  PIN io_logical_analyzer_packet[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 370.640 500.000 371.240 ;
    END
  END io_logical_analyzer_packet[67]
  PIN io_logical_analyzer_packet[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END io_logical_analyzer_packet[68]
  PIN io_logical_analyzer_packet[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END io_logical_analyzer_packet[69]
  PIN io_logical_analyzer_packet[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END io_logical_analyzer_packet[6]
  PIN io_logical_analyzer_packet[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_logical_analyzer_packet[70]
  PIN io_logical_analyzer_packet[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END io_logical_analyzer_packet[71]
  PIN io_logical_analyzer_packet[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END io_logical_analyzer_packet[72]
  PIN io_logical_analyzer_packet[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 796.000 435.070 800.000 ;
    END
  END io_logical_analyzer_packet[73]
  PIN io_logical_analyzer_packet[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.240 500.000 248.840 ;
    END
  END io_logical_analyzer_packet[74]
  PIN io_logical_analyzer_packet[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_logical_analyzer_packet[75]
  PIN io_logical_analyzer_packet[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 796.000 451.170 800.000 ;
    END
  END io_logical_analyzer_packet[76]
  PIN io_logical_analyzer_packet[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 796.000 278.670 800.000 ;
    END
  END io_logical_analyzer_packet[77]
  PIN io_logical_analyzer_packet[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_logical_analyzer_packet[78]
  PIN io_logical_analyzer_packet[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 796.000 299.370 800.000 ;
    END
  END io_logical_analyzer_packet[79]
  PIN io_logical_analyzer_packet[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 796.000 129.170 800.000 ;
    END
  END io_logical_analyzer_packet[7]
  PIN io_logical_analyzer_packet[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.040 500.000 459.640 ;
    END
  END io_logical_analyzer_packet[80]
  PIN io_logical_analyzer_packet[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 588.240 500.000 588.840 ;
    END
  END io_logical_analyzer_packet[81]
  PIN io_logical_analyzer_packet[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_logical_analyzer_packet[82]
  PIN io_logical_analyzer_packet[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 796.000 131.470 800.000 ;
    END
  END io_logical_analyzer_packet[83]
  PIN io_logical_analyzer_packet[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 520.240 500.000 520.840 ;
    END
  END io_logical_analyzer_packet[84]
  PIN io_logical_analyzer_packet[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END io_logical_analyzer_packet[85]
  PIN io_logical_analyzer_packet[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 796.000 126.870 800.000 ;
    END
  END io_logical_analyzer_packet[8]
  PIN io_logical_analyzer_packet[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 796.000 209.670 800.000 ;
    END
  END io_logical_analyzer_packet[9]
  PIN io_sram0_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END io_sram0_connections[0]
  PIN io_sram0_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 796.000 25.670 800.000 ;
    END
  END io_sram0_connections[10]
  PIN io_sram0_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END io_sram0_connections[11]
  PIN io_sram0_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 622.240 500.000 622.840 ;
    END
  END io_sram0_connections[12]
  PIN io_sram0_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END io_sram0_connections[13]
  PIN io_sram0_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 796.000 172.870 800.000 ;
    END
  END io_sram0_connections[14]
  PIN io_sram0_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END io_sram0_connections[15]
  PIN io_sram0_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 326.440 500.000 327.040 ;
    END
  END io_sram0_connections[16]
  PIN io_sram0_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END io_sram0_connections[17]
  PIN io_sram0_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END io_sram0_connections[18]
  PIN io_sram0_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END io_sram0_connections[19]
  PIN io_sram0_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 796.000 69.370 800.000 ;
    END
  END io_sram0_connections[1]
  PIN io_sram0_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 796.000 193.570 800.000 ;
    END
  END io_sram0_connections[20]
  PIN io_sram0_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END io_sram0_connections[21]
  PIN io_sram0_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_sram0_connections[22]
  PIN io_sram0_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 761.640 500.000 762.240 ;
    END
  END io_sram0_connections[23]
  PIN io_sram0_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_sram0_connections[24]
  PIN io_sram0_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END io_sram0_connections[25]
  PIN io_sram0_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END io_sram0_connections[26]
  PIN io_sram0_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END io_sram0_connections[27]
  PIN io_sram0_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 796.000 96.970 800.000 ;
    END
  END io_sram0_connections[28]
  PIN io_sram0_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 149.640 500.000 150.240 ;
    END
  END io_sram0_connections[29]
  PIN io_sram0_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 796.000 46.370 800.000 ;
    END
  END io_sram0_connections[2]
  PIN io_sram0_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END io_sram0_connections[30]
  PIN io_sram0_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_sram0_connections[31]
  PIN io_sram0_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_sram0_connections[32]
  PIN io_sram0_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 796.000 412.070 800.000 ;
    END
  END io_sram0_connections[33]
  PIN io_sram0_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 13.640 500.000 14.240 ;
    END
  END io_sram0_connections[34]
  PIN io_sram0_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 796.000 106.170 800.000 ;
    END
  END io_sram0_connections[35]
  PIN io_sram0_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 796.000 320.070 800.000 ;
    END
  END io_sram0_connections[36]
  PIN io_sram0_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 796.000 474.170 800.000 ;
    END
  END io_sram0_connections[37]
  PIN io_sram0_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 796.000 99.270 800.000 ;
    END
  END io_sram0_connections[38]
  PIN io_sram0_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 425.040 500.000 425.640 ;
    END
  END io_sram0_connections[39]
  PIN io_sram0_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END io_sram0_connections[3]
  PIN io_sram0_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 796.000 207.370 800.000 ;
    END
  END io_sram0_connections[40]
  PIN io_sram0_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_sram0_connections[41]
  PIN io_sram0_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 796.000 205.070 800.000 ;
    END
  END io_sram0_connections[42]
  PIN io_sram0_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 796.000 301.670 800.000 ;
    END
  END io_sram0_connections[43]
  PIN io_sram0_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.240 500.000 163.840 ;
    END
  END io_sram0_connections[44]
  PIN io_sram0_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END io_sram0_connections[45]
  PIN io_sram0_connections[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 710.640 500.000 711.240 ;
    END
  END io_sram0_connections[46]
  PIN io_sram0_connections[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 173.440 500.000 174.040 ;
    END
  END io_sram0_connections[47]
  PIN io_sram0_connections[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.840 500.000 398.440 ;
    END
  END io_sram0_connections[48]
  PIN io_sram0_connections[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END io_sram0_connections[49]
  PIN io_sram0_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 669.840 500.000 670.440 ;
    END
  END io_sram0_connections[4]
  PIN io_sram0_connections[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END io_sram0_connections[50]
  PIN io_sram0_connections[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END io_sram0_connections[51]
  PIN io_sram0_connections[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END io_sram0_connections[52]
  PIN io_sram0_connections[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END io_sram0_connections[53]
  PIN io_sram0_connections[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 765.040 500.000 765.640 ;
    END
  END io_sram0_connections[54]
  PIN io_sram0_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 122.440 500.000 123.040 ;
    END
  END io_sram0_connections[5]
  PIN io_sram0_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END io_sram0_connections[6]
  PIN io_sram0_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 796.000 359.170 800.000 ;
    END
  END io_sram0_connections[7]
  PIN io_sram0_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END io_sram0_connections[8]
  PIN io_sram0_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END io_sram0_connections[9]
  PIN io_sram0_r0_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 574.640 500.000 575.240 ;
    END
  END io_sram0_r0_in[0]
  PIN io_sram0_r0_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END io_sram0_r0_in[10]
  PIN io_sram0_r0_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 796.000 156.770 800.000 ;
    END
  END io_sram0_r0_in[11]
  PIN io_sram0_r0_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END io_sram0_r0_in[12]
  PIN io_sram0_r0_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 462.440 500.000 463.040 ;
    END
  END io_sram0_r0_in[13]
  PIN io_sram0_r0_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 81.640 500.000 82.240 ;
    END
  END io_sram0_r0_in[14]
  PIN io_sram0_r0_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_sram0_r0_in[15]
  PIN io_sram0_r0_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END io_sram0_r0_in[16]
  PIN io_sram0_r0_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 796.000 41.770 800.000 ;
    END
  END io_sram0_r0_in[17]
  PIN io_sram0_r0_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 796.000 416.670 800.000 ;
    END
  END io_sram0_r0_in[18]
  PIN io_sram0_r0_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 639.240 500.000 639.840 ;
    END
  END io_sram0_r0_in[19]
  PIN io_sram0_r0_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 788.840 500.000 789.440 ;
    END
  END io_sram0_r0_in[1]
  PIN io_sram0_r0_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 796.000 379.870 800.000 ;
    END
  END io_sram0_r0_in[20]
  PIN io_sram0_r0_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 796.000 347.670 800.000 ;
    END
  END io_sram0_r0_in[21]
  PIN io_sram0_r0_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END io_sram0_r0_in[22]
  PIN io_sram0_r0_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 796.000 285.570 800.000 ;
    END
  END io_sram0_r0_in[23]
  PIN io_sram0_r0_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END io_sram0_r0_in[24]
  PIN io_sram0_r0_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_sram0_r0_in[25]
  PIN io_sram0_r0_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_sram0_r0_in[26]
  PIN io_sram0_r0_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 796.000 487.970 800.000 ;
    END
  END io_sram0_r0_in[27]
  PIN io_sram0_r0_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END io_sram0_r0_in[28]
  PIN io_sram0_r0_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 374.040 500.000 374.640 ;
    END
  END io_sram0_r0_in[29]
  PIN io_sram0_r0_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END io_sram0_r0_in[2]
  PIN io_sram0_r0_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 796.000 161.370 800.000 ;
    END
  END io_sram0_r0_in[30]
  PIN io_sram0_r0_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 796.000 437.370 800.000 ;
    END
  END io_sram0_r0_in[31]
  PIN io_sram0_r0_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END io_sram0_r0_in[3]
  PIN io_sram0_r0_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 489.640 500.000 490.240 ;
    END
  END io_sram0_r0_in[4]
  PIN io_sram0_r0_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END io_sram0_r0_in[5]
  PIN io_sram0_r0_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_sram0_r0_in[6]
  PIN io_sram0_r0_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 792.240 500.000 792.840 ;
    END
  END io_sram0_r0_in[7]
  PIN io_sram0_r0_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 530.440 500.000 531.040 ;
    END
  END io_sram0_r0_in[8]
  PIN io_sram0_r0_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_sram0_r0_in[9]
  PIN io_sram0_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 796.000 469.570 800.000 ;
    END
  END io_sram0_rw_in[0]
  PIN io_sram0_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 782.040 500.000 782.640 ;
    END
  END io_sram0_rw_in[10]
  PIN io_sram0_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END io_sram0_rw_in[11]
  PIN io_sram0_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END io_sram0_rw_in[12]
  PIN io_sram0_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END io_sram0_rw_in[13]
  PIN io_sram0_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END io_sram0_rw_in[14]
  PIN io_sram0_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_sram0_rw_in[15]
  PIN io_sram0_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 796.000 14.170 800.000 ;
    END
  END io_sram0_rw_in[16]
  PIN io_sram0_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.840 500.000 347.440 ;
    END
  END io_sram0_rw_in[17]
  PIN io_sram0_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_sram0_rw_in[18]
  PIN io_sram0_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 673.240 500.000 673.840 ;
    END
  END io_sram0_rw_in[19]
  PIN io_sram0_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END io_sram0_rw_in[1]
  PIN io_sram0_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 796.000 60.170 800.000 ;
    END
  END io_sram0_rw_in[20]
  PIN io_sram0_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END io_sram0_rw_in[21]
  PIN io_sram0_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END io_sram0_rw_in[22]
  PIN io_sram0_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END io_sram0_rw_in[23]
  PIN io_sram0_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 207.440 500.000 208.040 ;
    END
  END io_sram0_rw_in[24]
  PIN io_sram0_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 796.000 113.070 800.000 ;
    END
  END io_sram0_rw_in[25]
  PIN io_sram0_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END io_sram0_rw_in[26]
  PIN io_sram0_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 796.000 322.370 800.000 ;
    END
  END io_sram0_rw_in[27]
  PIN io_sram0_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END io_sram0_rw_in[28]
  PIN io_sram0_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END io_sram0_rw_in[29]
  PIN io_sram0_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 445.440 500.000 446.040 ;
    END
  END io_sram0_rw_in[2]
  PIN io_sram0_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 796.000 230.370 800.000 ;
    END
  END io_sram0_rw_in[30]
  PIN io_sram0_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 748.040 500.000 748.640 ;
    END
  END io_sram0_rw_in[31]
  PIN io_sram0_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 796.000 152.170 800.000 ;
    END
  END io_sram0_rw_in[3]
  PIN io_sram0_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 796.000 345.370 800.000 ;
    END
  END io_sram0_rw_in[4]
  PIN io_sram0_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 758.240 500.000 758.840 ;
    END
  END io_sram0_rw_in[5]
  PIN io_sram0_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END io_sram0_rw_in[6]
  PIN io_sram0_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END io_sram0_rw_in[7]
  PIN io_sram0_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 612.040 500.000 612.640 ;
    END
  END io_sram0_rw_in[8]
  PIN io_sram0_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END io_sram0_rw_in[9]
  PIN io_sram1_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_sram1_connections[0]
  PIN io_sram1_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END io_sram1_connections[10]
  PIN io_sram1_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END io_sram1_connections[11]
  PIN io_sram1_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_sram1_connections[12]
  PIN io_sram1_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END io_sram1_connections[13]
  PIN io_sram1_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 632.440 500.000 633.040 ;
    END
  END io_sram1_connections[14]
  PIN io_sram1_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END io_sram1_connections[15]
  PIN io_sram1_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 547.440 500.000 548.040 ;
    END
  END io_sram1_connections[16]
  PIN io_sram1_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END io_sram1_connections[17]
  PIN io_sram1_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END io_sram1_connections[18]
  PIN io_sram1_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END io_sram1_connections[19]
  PIN io_sram1_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END io_sram1_connections[1]
  PIN io_sram1_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_sram1_connections[20]
  PIN io_sram1_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 741.240 500.000 741.840 ;
    END
  END io_sram1_connections[21]
  PIN io_sram1_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 796.000 239.570 800.000 ;
    END
  END io_sram1_connections[22]
  PIN io_sram1_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END io_sram1_connections[23]
  PIN io_sram1_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END io_sram1_connections[24]
  PIN io_sram1_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END io_sram1_connections[25]
  PIN io_sram1_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_sram1_connections[26]
  PIN io_sram1_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 796.000 409.770 800.000 ;
    END
  END io_sram1_connections[27]
  PIN io_sram1_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 796.000 115.370 800.000 ;
    END
  END io_sram1_connections[28]
  PIN io_sram1_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 796.000 356.870 800.000 ;
    END
  END io_sram1_connections[29]
  PIN io_sram1_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_sram1_connections[2]
  PIN io_sram1_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 578.040 500.000 578.640 ;
    END
  END io_sram1_connections[30]
  PIN io_sram1_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 697.040 500.000 697.640 ;
    END
  END io_sram1_connections[31]
  PIN io_sram1_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 796.000 117.670 800.000 ;
    END
  END io_sram1_connections[32]
  PIN io_sram1_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 796.000 124.570 800.000 ;
    END
  END io_sram1_connections[33]
  PIN io_sram1_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 796.000 395.970 800.000 ;
    END
  END io_sram1_connections[34]
  PIN io_sram1_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 796.000 382.170 800.000 ;
    END
  END io_sram1_connections[35]
  PIN io_sram1_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_sram1_connections[36]
  PIN io_sram1_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END io_sram1_connections[37]
  PIN io_sram1_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END io_sram1_connections[38]
  PIN io_sram1_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 796.000 253.370 800.000 ;
    END
  END io_sram1_connections[39]
  PIN io_sram1_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_sram1_connections[3]
  PIN io_sram1_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END io_sram1_connections[40]
  PIN io_sram1_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END io_sram1_connections[41]
  PIN io_sram1_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END io_sram1_connections[42]
  PIN io_sram1_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 796.000 7.270 800.000 ;
    END
  END io_sram1_connections[43]
  PIN io_sram1_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 796.000 241.870 800.000 ;
    END
  END io_sram1_connections[44]
  PIN io_sram1_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_sram1_connections[45]
  PIN io_sram1_connections[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END io_sram1_connections[46]
  PIN io_sram1_connections[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.040 500.000 170.640 ;
    END
  END io_sram1_connections[47]
  PIN io_sram1_connections[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 796.000 170.570 800.000 ;
    END
  END io_sram1_connections[48]
  PIN io_sram1_connections[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END io_sram1_connections[49]
  PIN io_sram1_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END io_sram1_connections[4]
  PIN io_sram1_connections[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 796.000 430.470 800.000 ;
    END
  END io_sram1_connections[50]
  PIN io_sram1_connections[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END io_sram1_connections[51]
  PIN io_sram1_connections[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_sram1_connections[52]
  PIN io_sram1_connections[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END io_sram1_connections[53]
  PIN io_sram1_connections[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 618.840 500.000 619.440 ;
    END
  END io_sram1_connections[54]
  PIN io_sram1_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 309.440 500.000 310.040 ;
    END
  END io_sram1_connections[5]
  PIN io_sram1_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_sram1_connections[6]
  PIN io_sram1_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 796.000 441.970 800.000 ;
    END
  END io_sram1_connections[7]
  PIN io_sram1_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 391.040 500.000 391.640 ;
    END
  END io_sram1_connections[8]
  PIN io_sram1_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END io_sram1_connections[9]
  PIN io_sram1_ro_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END io_sram1_ro_in[0]
  PIN io_sram1_ro_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_sram1_ro_in[10]
  PIN io_sram1_ro_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END io_sram1_ro_in[11]
  PIN io_sram1_ro_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END io_sram1_ro_in[12]
  PIN io_sram1_ro_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_sram1_ro_in[13]
  PIN io_sram1_ro_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 796.000 4.970 800.000 ;
    END
  END io_sram1_ro_in[14]
  PIN io_sram1_ro_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 796.000 11.870 800.000 ;
    END
  END io_sram1_ro_in[15]
  PIN io_sram1_ro_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 796.000 361.470 800.000 ;
    END
  END io_sram1_ro_in[16]
  PIN io_sram1_ro_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END io_sram1_ro_in[17]
  PIN io_sram1_ro_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 190.440 500.000 191.040 ;
    END
  END io_sram1_ro_in[18]
  PIN io_sram1_ro_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END io_sram1_ro_in[19]
  PIN io_sram1_ro_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END io_sram1_ro_in[1]
  PIN io_sram1_ro_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 469.240 500.000 469.840 ;
    END
  END io_sram1_ro_in[20]
  PIN io_sram1_ro_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END io_sram1_ro_in[21]
  PIN io_sram1_ro_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 796.000 218.870 800.000 ;
    END
  END io_sram1_ro_in[22]
  PIN io_sram1_ro_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END io_sram1_ro_in[23]
  PIN io_sram1_ro_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END io_sram1_ro_in[24]
  PIN io_sram1_ro_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END io_sram1_ro_in[25]
  PIN io_sram1_ro_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END io_sram1_ro_in[26]
  PIN io_sram1_ro_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END io_sram1_ro_in[27]
  PIN io_sram1_ro_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END io_sram1_ro_in[28]
  PIN io_sram1_ro_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END io_sram1_ro_in[29]
  PIN io_sram1_ro_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.240 500.000 27.840 ;
    END
  END io_sram1_ro_in[2]
  PIN io_sram1_ro_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END io_sram1_ro_in[30]
  PIN io_sram1_ro_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_sram1_ro_in[31]
  PIN io_sram1_ro_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_sram1_ro_in[3]
  PIN io_sram1_ro_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 796.000 53.270 800.000 ;
    END
  END io_sram1_ro_in[4]
  PIN io_sram1_ro_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END io_sram1_ro_in[5]
  PIN io_sram1_ro_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.040 500.000 204.640 ;
    END
  END io_sram1_ro_in[6]
  PIN io_sram1_ro_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END io_sram1_ro_in[7]
  PIN io_sram1_ro_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 438.640 500.000 439.240 ;
    END
  END io_sram1_ro_in[8]
  PIN io_sram1_ro_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 796.000 64.770 800.000 ;
    END
  END io_sram1_ro_in[9]
  PIN io_sram1_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END io_sram1_rw_in[0]
  PIN io_sram1_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_sram1_rw_in[10]
  PIN io_sram1_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 796.000 471.870 800.000 ;
    END
  END io_sram1_rw_in[11]
  PIN io_sram1_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END io_sram1_rw_in[12]
  PIN io_sram1_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 533.840 500.000 534.440 ;
    END
  END io_sram1_rw_in[13]
  PIN io_sram1_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END io_sram1_rw_in[14]
  PIN io_sram1_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END io_sram1_rw_in[15]
  PIN io_sram1_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 796.000 76.270 800.000 ;
    END
  END io_sram1_rw_in[16]
  PIN io_sram1_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END io_sram1_rw_in[17]
  PIN io_sram1_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 129.240 500.000 129.840 ;
    END
  END io_sram1_rw_in[18]
  PIN io_sram1_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 37.440 500.000 38.040 ;
    END
  END io_sram1_rw_in[19]
  PIN io_sram1_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 751.440 500.000 752.040 ;
    END
  END io_sram1_rw_in[1]
  PIN io_sram1_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 54.440 500.000 55.040 ;
    END
  END io_sram1_rw_in[20]
  PIN io_sram1_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 754.840 500.000 755.440 ;
    END
  END io_sram1_rw_in[21]
  PIN io_sram1_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_sram1_rw_in[22]
  PIN io_sram1_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 796.000 221.170 800.000 ;
    END
  END io_sram1_rw_in[23]
  PIN io_sram1_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 796.000 405.170 800.000 ;
    END
  END io_sram1_rw_in[24]
  PIN io_sram1_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 394.440 500.000 395.040 ;
    END
  END io_sram1_rw_in[25]
  PIN io_sram1_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END io_sram1_rw_in[26]
  PIN io_sram1_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_sram1_rw_in[27]
  PIN io_sram1_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_sram1_rw_in[28]
  PIN io_sram1_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END io_sram1_rw_in[29]
  PIN io_sram1_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END io_sram1_rw_in[2]
  PIN io_sram1_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END io_sram1_rw_in[30]
  PIN io_sram1_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 796.000 94.670 800.000 ;
    END
  END io_sram1_rw_in[31]
  PIN io_sram1_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 734.440 500.000 735.040 ;
    END
  END io_sram1_rw_in[3]
  PIN io_sram1_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 455.640 500.000 456.240 ;
    END
  END io_sram1_rw_in[4]
  PIN io_sram1_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.840 500.000 279.440 ;
    END
  END io_sram1_rw_in[5]
  PIN io_sram1_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 47.640 500.000 48.240 ;
    END
  END io_sram1_rw_in[6]
  PIN io_sram1_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 796.000 494.870 800.000 ;
    END
  END io_sram1_rw_in[7]
  PIN io_sram1_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 796.000 44.070 800.000 ;
    END
  END io_sram1_rw_in[8]
  PIN io_sram1_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END io_sram1_rw_in[9]
  PIN io_sram2_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END io_sram2_connections[0]
  PIN io_sram2_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 796.000 30.270 800.000 ;
    END
  END io_sram2_connections[10]
  PIN io_sram2_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.240 500.000 146.840 ;
    END
  END io_sram2_connections[11]
  PIN io_sram2_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 503.240 500.000 503.840 ;
    END
  END io_sram2_connections[12]
  PIN io_sram2_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 796.000 165.970 800.000 ;
    END
  END io_sram2_connections[13]
  PIN io_sram2_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_sram2_connections[14]
  PIN io_sram2_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END io_sram2_connections[15]
  PIN io_sram2_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 796.000 336.170 800.000 ;
    END
  END io_sram2_connections[16]
  PIN io_sram2_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 656.240 500.000 656.840 ;
    END
  END io_sram2_connections[17]
  PIN io_sram2_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END io_sram2_connections[18]
  PIN io_sram2_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END io_sram2_connections[19]
  PIN io_sram2_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END io_sram2_connections[1]
  PIN io_sram2_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 796.000 418.970 800.000 ;
    END
  END io_sram2_connections[20]
  PIN io_sram2_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 796.000 119.970 800.000 ;
    END
  END io_sram2_connections[21]
  PIN io_sram2_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_sram2_connections[22]
  PIN io_sram2_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.840 500.000 313.440 ;
    END
  END io_sram2_connections[23]
  PIN io_sram2_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_sram2_connections[24]
  PIN io_sram2_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_sram2_connections[25]
  PIN io_sram2_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END io_sram2_connections[26]
  PIN io_sram2_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END io_sram2_connections[27]
  PIN io_sram2_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 796.000 384.470 800.000 ;
    END
  END io_sram2_connections[28]
  PIN io_sram2_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END io_sram2_connections[29]
  PIN io_sram2_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_sram2_connections[2]
  PIN io_sram2_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 796.000 103.870 800.000 ;
    END
  END io_sram2_connections[30]
  PIN io_sram2_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io_sram2_connections[31]
  PIN io_sram2_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 796.000 110.770 800.000 ;
    END
  END io_sram2_connections[32]
  PIN io_sram2_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END io_sram2_connections[33]
  PIN io_sram2_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END io_sram2_connections[34]
  PIN io_sram2_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 796.000 402.870 800.000 ;
    END
  END io_sram2_connections[35]
  PIN io_sram2_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END io_sram2_connections[36]
  PIN io_sram2_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 796.000 87.770 800.000 ;
    END
  END io_sram2_connections[37]
  PIN io_sram2_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 796.000 21.070 800.000 ;
    END
  END io_sram2_connections[38]
  PIN io_sram2_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END io_sram2_connections[39]
  PIN io_sram2_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END io_sram2_connections[3]
  PIN io_sram2_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_sram2_connections[40]
  PIN io_sram2_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 796.000 48.670 800.000 ;
    END
  END io_sram2_connections[41]
  PIN io_sram2_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 796.000 414.370 800.000 ;
    END
  END io_sram2_connections[42]
  PIN io_sram2_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END io_sram2_connections[43]
  PIN io_sram2_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io_sram2_connections[44]
  PIN io_sram2_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 506.640 500.000 507.240 ;
    END
  END io_sram2_connections[45]
  PIN io_sram2_connections[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END io_sram2_connections[46]
  PIN io_sram2_connections[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END io_sram2_connections[47]
  PIN io_sram2_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.840 500.000 296.440 ;
    END
  END io_sram2_connections[4]
  PIN io_sram2_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 10.240 500.000 10.840 ;
    END
  END io_sram2_connections[5]
  PIN io_sram2_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END io_sram2_connections[6]
  PIN io_sram2_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END io_sram2_connections[7]
  PIN io_sram2_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END io_sram2_connections[8]
  PIN io_sram2_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_sram2_connections[9]
  PIN io_sram2_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 350.240 500.000 350.840 ;
    END
  END io_sram2_rw_in[0]
  PIN io_sram2_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.240 500.000 282.840 ;
    END
  END io_sram2_rw_in[10]
  PIN io_sram2_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 567.840 500.000 568.440 ;
    END
  END io_sram2_rw_in[11]
  PIN io_sram2_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 292.440 500.000 293.040 ;
    END
  END io_sram2_rw_in[12]
  PIN io_sram2_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END io_sram2_rw_in[13]
  PIN io_sram2_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 796.000 324.670 800.000 ;
    END
  END io_sram2_rw_in[14]
  PIN io_sram2_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END io_sram2_rw_in[15]
  PIN io_sram2_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END io_sram2_rw_in[16]
  PIN io_sram2_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 796.000 264.870 800.000 ;
    END
  END io_sram2_rw_in[17]
  PIN io_sram2_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.240 500.000 214.840 ;
    END
  END io_sram2_rw_in[18]
  PIN io_sram2_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END io_sram2_rw_in[19]
  PIN io_sram2_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 771.840 500.000 772.440 ;
    END
  END io_sram2_rw_in[1]
  PIN io_sram2_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 796.000 444.270 800.000 ;
    END
  END io_sram2_rw_in[20]
  PIN io_sram2_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 591.640 500.000 592.240 ;
    END
  END io_sram2_rw_in[21]
  PIN io_sram2_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END io_sram2_rw_in[22]
  PIN io_sram2_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_sram2_rw_in[23]
  PIN io_sram2_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 796.000 310.870 800.000 ;
    END
  END io_sram2_rw_in[24]
  PIN io_sram2_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END io_sram2_rw_in[25]
  PIN io_sram2_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END io_sram2_rw_in[26]
  PIN io_sram2_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END io_sram2_rw_in[27]
  PIN io_sram2_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_sram2_rw_in[28]
  PIN io_sram2_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END io_sram2_rw_in[29]
  PIN io_sram2_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END io_sram2_rw_in[2]
  PIN io_sram2_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 778.640 500.000 779.240 ;
    END
  END io_sram2_rw_in[30]
  PIN io_sram2_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 115.640 500.000 116.240 ;
    END
  END io_sram2_rw_in[31]
  PIN io_sram2_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END io_sram2_rw_in[3]
  PIN io_sram2_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END io_sram2_rw_in[4]
  PIN io_sram2_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END io_sram2_rw_in[5]
  PIN io_sram2_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END io_sram2_rw_in[6]
  PIN io_sram2_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_sram2_rw_in[7]
  PIN io_sram2_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 796.000 198.170 800.000 ;
    END
  END io_sram2_rw_in[8]
  PIN io_sram2_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_sram2_rw_in[9]
  PIN io_sram3_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END io_sram3_connections[0]
  PIN io_sram3_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END io_sram3_connections[10]
  PIN io_sram3_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io_sram3_connections[11]
  PIN io_sram3_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 796.000 232.670 800.000 ;
    END
  END io_sram3_connections[12]
  PIN io_sram3_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END io_sram3_connections[13]
  PIN io_sram3_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_sram3_connections[14]
  PIN io_sram3_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 479.440 500.000 480.040 ;
    END
  END io_sram3_connections[15]
  PIN io_sram3_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 796.000 460.370 800.000 ;
    END
  END io_sram3_connections[16]
  PIN io_sram3_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END io_sram3_connections[17]
  PIN io_sram3_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END io_sram3_connections[18]
  PIN io_sram3_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 796.000 78.570 800.000 ;
    END
  END io_sram3_connections[19]
  PIN io_sram3_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 796.000 271.770 800.000 ;
    END
  END io_sram3_connections[1]
  PIN io_sram3_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.240 500.000 61.840 ;
    END
  END io_sram3_connections[20]
  PIN io_sram3_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.840 500.000 194.440 ;
    END
  END io_sram3_connections[21]
  PIN io_sram3_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_sram3_connections[22]
  PIN io_sram3_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 796.000 188.970 800.000 ;
    END
  END io_sram3_connections[23]
  PIN io_sram3_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END io_sram3_connections[24]
  PIN io_sram3_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END io_sram3_connections[25]
  PIN io_sram3_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_sram3_connections[26]
  PIN io_sram3_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 768.440 500.000 769.040 ;
    END
  END io_sram3_connections[27]
  PIN io_sram3_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 663.040 500.000 663.640 ;
    END
  END io_sram3_connections[28]
  PIN io_sram3_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END io_sram3_connections[29]
  PIN io_sram3_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END io_sram3_connections[2]
  PIN io_sram3_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_sram3_connections[30]
  PIN io_sram3_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END io_sram3_connections[31]
  PIN io_sram3_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END io_sram3_connections[32]
  PIN io_sram3_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END io_sram3_connections[33]
  PIN io_sram3_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_sram3_connections[34]
  PIN io_sram3_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END io_sram3_connections[35]
  PIN io_sram3_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END io_sram3_connections[36]
  PIN io_sram3_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 737.840 500.000 738.440 ;
    END
  END io_sram3_connections[37]
  PIN io_sram3_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END io_sram3_connections[38]
  PIN io_sram3_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 635.840 500.000 636.440 ;
    END
  END io_sram3_connections[39]
  PIN io_sram3_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 796.000 400.570 800.000 ;
    END
  END io_sram3_connections[3]
  PIN io_sram3_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_sram3_connections[40]
  PIN io_sram3_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END io_sram3_connections[41]
  PIN io_sram3_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 796.000 478.770 800.000 ;
    END
  END io_sram3_connections[42]
  PIN io_sram3_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END io_sram3_connections[43]
  PIN io_sram3_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 796.000 317.770 800.000 ;
    END
  END io_sram3_connections[44]
  PIN io_sram3_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END io_sram3_connections[45]
  PIN io_sram3_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 796.000 262.570 800.000 ;
    END
  END io_sram3_connections[4]
  PIN io_sram3_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 78.240 500.000 78.840 ;
    END
  END io_sram3_connections[5]
  PIN io_sram3_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END io_sram3_connections[6]
  PIN io_sram3_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_sram3_connections[7]
  PIN io_sram3_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 608.640 500.000 609.240 ;
    END
  END io_sram3_connections[8]
  PIN io_sram3_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 796.000 159.070 800.000 ;
    END
  END io_sram3_connections[9]
  PIN io_sram3_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END io_sram3_rw_in[0]
  PIN io_sram3_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 796.000 133.770 800.000 ;
    END
  END io_sram3_rw_in[10]
  PIN io_sram3_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 183.640 500.000 184.240 ;
    END
  END io_sram3_rw_in[11]
  PIN io_sram3_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 540.640 500.000 541.240 ;
    END
  END io_sram3_rw_in[12]
  PIN io_sram3_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_sram3_rw_in[13]
  PIN io_sram3_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.840 500.000 415.440 ;
    END
  END io_sram3_rw_in[14]
  PIN io_sram3_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_sram3_rw_in[15]
  PIN io_sram3_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 323.040 500.000 323.640 ;
    END
  END io_sram3_rw_in[16]
  PIN io_sram3_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END io_sram3_rw_in[17]
  PIN io_sram3_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END io_sram3_rw_in[18]
  PIN io_sram3_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 690.240 500.000 690.840 ;
    END
  END io_sram3_rw_in[19]
  PIN io_sram3_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.840 500.000 449.440 ;
    END
  END io_sram3_rw_in[1]
  PIN io_sram3_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END io_sram3_rw_in[20]
  PIN io_sram3_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io_sram3_rw_in[21]
  PIN io_sram3_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END io_sram3_rw_in[22]
  PIN io_sram3_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END io_sram3_rw_in[23]
  PIN io_sram3_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 785.440 500.000 786.040 ;
    END
  END io_sram3_rw_in[24]
  PIN io_sram3_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END io_sram3_rw_in[25]
  PIN io_sram3_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END io_sram3_rw_in[26]
  PIN io_sram3_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END io_sram3_rw_in[27]
  PIN io_sram3_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 796.000 338.470 800.000 ;
    END
  END io_sram3_rw_in[28]
  PIN io_sram3_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END io_sram3_rw_in[29]
  PIN io_sram3_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 625.640 500.000 626.240 ;
    END
  END io_sram3_rw_in[2]
  PIN io_sram3_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 796.000 497.170 800.000 ;
    END
  END io_sram3_rw_in[30]
  PIN io_sram3_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END io_sram3_rw_in[31]
  PIN io_sram3_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END io_sram3_rw_in[3]
  PIN io_sram3_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 796.000 492.570 800.000 ;
    END
  END io_sram3_rw_in[4]
  PIN io_sram3_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END io_sram3_rw_in[5]
  PIN io_sram3_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END io_sram3_rw_in[6]
  PIN io_sram3_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END io_sram3_rw_in[7]
  PIN io_sram3_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 796.000 260.270 800.000 ;
    END
  END io_sram3_rw_in[8]
  PIN io_sram3_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 796.000 18.770 800.000 ;
    END
  END io_sram3_rw_in[9]
  PIN io_sram4_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 796.000 136.070 800.000 ;
    END
  END io_sram4_connections[0]
  PIN io_sram4_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 336.640 500.000 337.240 ;
    END
  END io_sram4_connections[10]
  PIN io_sram4_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END io_sram4_connections[11]
  PIN io_sram4_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END io_sram4_connections[12]
  PIN io_sram4_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 717.440 500.000 718.040 ;
    END
  END io_sram4_connections[13]
  PIN io_sram4_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_sram4_connections[14]
  PIN io_sram4_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 796.000 37.170 800.000 ;
    END
  END io_sram4_connections[15]
  PIN io_sram4_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END io_sram4_connections[16]
  PIN io_sram4_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END io_sram4_connections[17]
  PIN io_sram4_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_sram4_connections[18]
  PIN io_sram4_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_sram4_connections[19]
  PIN io_sram4_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END io_sram4_connections[1]
  PIN io_sram4_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 796.000 195.870 800.000 ;
    END
  END io_sram4_connections[20]
  PIN io_sram4_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END io_sram4_connections[21]
  PIN io_sram4_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 796.000 292.470 800.000 ;
    END
  END io_sram4_connections[22]
  PIN io_sram4_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 435.240 500.000 435.840 ;
    END
  END io_sram4_connections[23]
  PIN io_sram4_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 796.000 326.970 800.000 ;
    END
  END io_sram4_connections[24]
  PIN io_sram4_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 796.000 455.770 800.000 ;
    END
  END io_sram4_connections[25]
  PIN io_sram4_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_sram4_connections[26]
  PIN io_sram4_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 227.840 500.000 228.440 ;
    END
  END io_sram4_connections[27]
  PIN io_sram4_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END io_sram4_connections[28]
  PIN io_sram4_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END io_sram4_connections[29]
  PIN io_sram4_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END io_sram4_connections[2]
  PIN io_sram4_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END io_sram4_connections[30]
  PIN io_sram4_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END io_sram4_connections[31]
  PIN io_sram4_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 796.000 140.670 800.000 ;
    END
  END io_sram4_connections[32]
  PIN io_sram4_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 795.640 500.000 796.240 ;
    END
  END io_sram4_connections[33]
  PIN io_sram4_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END io_sram4_connections[34]
  PIN io_sram4_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END io_sram4_connections[35]
  PIN io_sram4_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 796.000 175.170 800.000 ;
    END
  END io_sram4_connections[36]
  PIN io_sram4_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_sram4_connections[37]
  PIN io_sram4_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.840 500.000 364.440 ;
    END
  END io_sram4_connections[38]
  PIN io_sram4_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END io_sram4_connections[39]
  PIN io_sram4_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END io_sram4_connections[3]
  PIN io_sram4_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 796.000 71.670 800.000 ;
    END
  END io_sram4_connections[40]
  PIN io_sram4_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END io_sram4_connections[41]
  PIN io_sram4_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 796.000 186.670 800.000 ;
    END
  END io_sram4_connections[42]
  PIN io_sram4_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 659.640 500.000 660.240 ;
    END
  END io_sram4_connections[43]
  PIN io_sram4_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 796.000 90.070 800.000 ;
    END
  END io_sram4_connections[44]
  PIN io_sram4_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END io_sram4_connections[45]
  PIN io_sram4_connections[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_sram4_connections[46]
  PIN io_sram4_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 493.040 500.000 493.640 ;
    END
  END io_sram4_connections[4]
  PIN io_sram4_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END io_sram4_connections[5]
  PIN io_sram4_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END io_sram4_connections[6]
  PIN io_sram4_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END io_sram4_connections[7]
  PIN io_sram4_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.040 500.000 17.640 ;
    END
  END io_sram4_connections[8]
  PIN io_sram4_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.040 500.000 119.640 ;
    END
  END io_sram4_connections[9]
  PIN io_sram4_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 796.000 421.270 800.000 ;
    END
  END io_sram4_rw_in[0]
  PIN io_sram4_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 796.000 80.870 800.000 ;
    END
  END io_sram4_rw_in[10]
  PIN io_sram4_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_sram4_rw_in[11]
  PIN io_sram4_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END io_sram4_rw_in[12]
  PIN io_sram4_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 796.000 386.770 800.000 ;
    END
  END io_sram4_rw_in[13]
  PIN io_sram4_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 680.040 500.000 680.640 ;
    END
  END io_sram4_rw_in[14]
  PIN io_sram4_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 796.000 228.070 800.000 ;
    END
  END io_sram4_rw_in[15]
  PIN io_sram4_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END io_sram4_rw_in[16]
  PIN io_sram4_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END io_sram4_rw_in[17]
  PIN io_sram4_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END io_sram4_rw_in[18]
  PIN io_sram4_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 700.440 500.000 701.040 ;
    END
  END io_sram4_rw_in[19]
  PIN io_sram4_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 796.000 237.270 800.000 ;
    END
  END io_sram4_rw_in[1]
  PIN io_sram4_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_sram4_rw_in[20]
  PIN io_sram4_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END io_sram4_rw_in[21]
  PIN io_sram4_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END io_sram4_rw_in[22]
  PIN io_sram4_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END io_sram4_rw_in[23]
  PIN io_sram4_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END io_sram4_rw_in[24]
  PIN io_sram4_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 796.000 182.070 800.000 ;
    END
  END io_sram4_rw_in[25]
  PIN io_sram4_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_sram4_rw_in[26]
  PIN io_sram4_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 601.840 500.000 602.440 ;
    END
  END io_sram4_rw_in[27]
  PIN io_sram4_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 796.000 276.370 800.000 ;
    END
  END io_sram4_rw_in[28]
  PIN io_sram4_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 200.640 500.000 201.240 ;
    END
  END io_sram4_rw_in[29]
  PIN io_sram4_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END io_sram4_rw_in[2]
  PIN io_sram4_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END io_sram4_rw_in[30]
  PIN io_sram4_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 796.000 464.970 800.000 ;
    END
  END io_sram4_rw_in[31]
  PIN io_sram4_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 796.000 375.270 800.000 ;
    END
  END io_sram4_rw_in[3]
  PIN io_sram4_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END io_sram4_rw_in[4]
  PIN io_sram4_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 796.000 290.170 800.000 ;
    END
  END io_sram4_rw_in[5]
  PIN io_sram4_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_sram4_rw_in[6]
  PIN io_sram4_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END io_sram4_rw_in[7]
  PIN io_sram4_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 649.440 500.000 650.040 ;
    END
  END io_sram4_rw_in[8]
  PIN io_sram4_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 561.040 500.000 561.640 ;
    END
  END io_sram4_rw_in[9]
  PIN io_sram5_connections[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END io_sram5_connections[0]
  PIN io_sram5_connections[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 796.000 340.770 800.000 ;
    END
  END io_sram5_connections[10]
  PIN io_sram5_connections[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 796.000 142.970 800.000 ;
    END
  END io_sram5_connections[11]
  PIN io_sram5_connections[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_sram5_connections[12]
  PIN io_sram5_connections[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 796.000 398.270 800.000 ;
    END
  END io_sram5_connections[13]
  PIN io_sram5_connections[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 796.000 145.270 800.000 ;
    END
  END io_sram5_connections[14]
  PIN io_sram5_connections[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 796.000 349.970 800.000 ;
    END
  END io_sram5_connections[15]
  PIN io_sram5_connections[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 720.840 500.000 721.440 ;
    END
  END io_sram5_connections[16]
  PIN io_sram5_connections[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_sram5_connections[17]
  PIN io_sram5_connections[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END io_sram5_connections[18]
  PIN io_sram5_connections[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 299.240 500.000 299.840 ;
    END
  END io_sram5_connections[19]
  PIN io_sram5_connections[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 302.640 500.000 303.240 ;
    END
  END io_sram5_connections[1]
  PIN io_sram5_connections[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_sram5_connections[20]
  PIN io_sram5_connections[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 796.000 313.170 800.000 ;
    END
  END io_sram5_connections[21]
  PIN io_sram5_connections[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END io_sram5_connections[22]
  PIN io_sram5_connections[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_sram5_connections[23]
  PIN io_sram5_connections[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END io_sram5_connections[24]
  PIN io_sram5_connections[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 744.640 500.000 745.240 ;
    END
  END io_sram5_connections[25]
  PIN io_sram5_connections[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_sram5_connections[26]
  PIN io_sram5_connections[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 652.840 500.000 653.440 ;
    END
  END io_sram5_connections[27]
  PIN io_sram5_connections[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END io_sram5_connections[28]
  PIN io_sram5_connections[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END io_sram5_connections[29]
  PIN io_sram5_connections[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.840 500.000 432.440 ;
    END
  END io_sram5_connections[2]
  PIN io_sram5_connections[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END io_sram5_connections[30]
  PIN io_sram5_connections[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END io_sram5_connections[31]
  PIN io_sram5_connections[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 796.000 9.570 800.000 ;
    END
  END io_sram5_connections[32]
  PIN io_sram5_connections[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_sram5_connections[33]
  PIN io_sram5_connections[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END io_sram5_connections[34]
  PIN io_sram5_connections[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END io_sram5_connections[35]
  PIN io_sram5_connections[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 6.840 500.000 7.440 ;
    END
  END io_sram5_connections[36]
  PIN io_sram5_connections[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 796.000 448.870 800.000 ;
    END
  END io_sram5_connections[37]
  PIN io_sram5_connections[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END io_sram5_connections[38]
  PIN io_sram5_connections[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 268.640 500.000 269.240 ;
    END
  END io_sram5_connections[39]
  PIN io_sram5_connections[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 796.000 149.870 800.000 ;
    END
  END io_sram5_connections[3]
  PIN io_sram5_connections[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END io_sram5_connections[40]
  PIN io_sram5_connections[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_sram5_connections[41]
  PIN io_sram5_connections[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END io_sram5_connections[42]
  PIN io_sram5_connections[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 595.040 500.000 595.640 ;
    END
  END io_sram5_connections[43]
  PIN io_sram5_connections[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 796.000 329.270 800.000 ;
    END
  END io_sram5_connections[44]
  PIN io_sram5_connections[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END io_sram5_connections[45]
  PIN io_sram5_connections[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 550.840 500.000 551.440 ;
    END
  END io_sram5_connections[46]
  PIN io_sram5_connections[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_sram5_connections[47]
  PIN io_sram5_connections[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 683.440 500.000 684.040 ;
    END
  END io_sram5_connections[48]
  PIN io_sram5_connections[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END io_sram5_connections[49]
  PIN io_sram5_connections[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END io_sram5_connections[4]
  PIN io_sram5_connections[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 316.240 500.000 316.840 ;
    END
  END io_sram5_connections[50]
  PIN io_sram5_connections[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.240 500.000 367.840 ;
    END
  END io_sram5_connections[51]
  PIN io_sram5_connections[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END io_sram5_connections[52]
  PIN io_sram5_connections[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_sram5_connections[53]
  PIN io_sram5_connections[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_sram5_connections[54]
  PIN io_sram5_connections[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 499.840 500.000 500.440 ;
    END
  END io_sram5_connections[55]
  PIN io_sram5_connections[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END io_sram5_connections[56]
  PIN io_sram5_connections[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.840 500.000 143.440 ;
    END
  END io_sram5_connections[57]
  PIN io_sram5_connections[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 353.640 500.000 354.240 ;
    END
  END io_sram5_connections[58]
  PIN io_sram5_connections[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 571.240 500.000 571.840 ;
    END
  END io_sram5_connections[59]
  PIN io_sram5_connections[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END io_sram5_connections[5]
  PIN io_sram5_connections[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END io_sram5_connections[60]
  PIN io_sram5_connections[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 796.000 57.870 800.000 ;
    END
  END io_sram5_connections[61]
  PIN io_sram5_connections[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END io_sram5_connections[62]
  PIN io_sram5_connections[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_sram5_connections[63]
  PIN io_sram5_connections[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_sram5_connections[64]
  PIN io_sram5_connections[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END io_sram5_connections[65]
  PIN io_sram5_connections[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_sram5_connections[66]
  PIN io_sram5_connections[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 796.000 251.070 800.000 ;
    END
  END io_sram5_connections[67]
  PIN io_sram5_connections[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END io_sram5_connections[68]
  PIN io_sram5_connections[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_sram5_connections[69]
  PIN io_sram5_connections[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END io_sram5_connections[6]
  PIN io_sram5_connections[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END io_sram5_connections[70]
  PIN io_sram5_connections[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_sram5_connections[71]
  PIN io_sram5_connections[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 544.040 500.000 544.640 ;
    END
  END io_sram5_connections[72]
  PIN io_sram5_connections[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END io_sram5_connections[73]
  PIN io_sram5_connections[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.240 500.000 384.840 ;
    END
  END io_sram5_connections[74]
  PIN io_sram5_connections[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 796.000 368.370 800.000 ;
    END
  END io_sram5_connections[75]
  PIN io_sram5_connections[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END io_sram5_connections[76]
  PIN io_sram5_connections[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_sram5_connections[77]
  PIN io_sram5_connections[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.040 500.000 476.640 ;
    END
  END io_sram5_connections[78]
  PIN io_sram5_connections[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 796.000 108.470 800.000 ;
    END
  END io_sram5_connections[79]
  PIN io_sram5_connections[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 796.000 377.570 800.000 ;
    END
  END io_sram5_connections[7]
  PIN io_sram5_connections[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END io_sram5_connections[80]
  PIN io_sram5_connections[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 796.000 246.470 800.000 ;
    END
  END io_sram5_connections[81]
  PIN io_sram5_connections[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END io_sram5_connections[82]
  PIN io_sram5_connections[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END io_sram5_connections[8]
  PIN io_sram5_connections[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END io_sram5_connections[9]
  PIN io_sram5_rw_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_sram5_rw_in[0]
  PIN io_sram5_rw_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 796.000 255.670 800.000 ;
    END
  END io_sram5_rw_in[10]
  PIN io_sram5_rw_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_sram5_rw_in[11]
  PIN io_sram5_rw_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END io_sram5_rw_in[12]
  PIN io_sram5_rw_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 584.840 500.000 585.440 ;
    END
  END io_sram5_rw_in[13]
  PIN io_sram5_rw_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 796.000 211.970 800.000 ;
    END
  END io_sram5_rw_in[14]
  PIN io_sram5_rw_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_sram5_rw_in[15]
  PIN io_sram5_rw_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END io_sram5_rw_in[16]
  PIN io_sram5_rw_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_sram5_rw_in[17]
  PIN io_sram5_rw_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 472.640 500.000 473.240 ;
    END
  END io_sram5_rw_in[18]
  PIN io_sram5_rw_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END io_sram5_rw_in[19]
  PIN io_sram5_rw_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END io_sram5_rw_in[1]
  PIN io_sram5_rw_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END io_sram5_rw_in[20]
  PIN io_sram5_rw_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 796.000 283.270 800.000 ;
    END
  END io_sram5_rw_in[21]
  PIN io_sram5_rw_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 796.000 315.470 800.000 ;
    END
  END io_sram5_rw_in[22]
  PIN io_sram5_rw_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END io_sram5_rw_in[23]
  PIN io_sram5_rw_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END io_sram5_rw_in[24]
  PIN io_sram5_rw_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 796.000 34.870 800.000 ;
    END
  END io_sram5_rw_in[25]
  PIN io_sram5_rw_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END io_sram5_rw_in[26]
  PIN io_sram5_rw_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 796.000 372.970 800.000 ;
    END
  END io_sram5_rw_in[27]
  PIN io_sram5_rw_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_sram5_rw_in[28]
  PIN io_sram5_rw_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END io_sram5_rw_in[29]
  PIN io_sram5_rw_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END io_sram5_rw_in[2]
  PIN io_sram5_rw_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END io_sram5_rw_in[30]
  PIN io_sram5_rw_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END io_sram5_rw_in[31]
  PIN io_sram5_rw_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END io_sram5_rw_in[32]
  PIN io_sram5_rw_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.840 500.000 75.440 ;
    END
  END io_sram5_rw_in[33]
  PIN io_sram5_rw_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END io_sram5_rw_in[34]
  PIN io_sram5_rw_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 796.000 267.170 800.000 ;
    END
  END io_sram5_rw_in[35]
  PIN io_sram5_rw_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_sram5_rw_in[36]
  PIN io_sram5_rw_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END io_sram5_rw_in[37]
  PIN io_sram5_rw_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.240 500.000 231.840 ;
    END
  END io_sram5_rw_in[38]
  PIN io_sram5_rw_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_sram5_rw_in[39]
  PIN io_sram5_rw_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 796.000 467.270 800.000 ;
    END
  END io_sram5_rw_in[3]
  PIN io_sram5_rw_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 796.000 476.470 800.000 ;
    END
  END io_sram5_rw_in[40]
  PIN io_sram5_rw_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_sram5_rw_in[41]
  PIN io_sram5_rw_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END io_sram5_rw_in[42]
  PIN io_sram5_rw_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_sram5_rw_in[43]
  PIN io_sram5_rw_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_sram5_rw_in[44]
  PIN io_sram5_rw_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END io_sram5_rw_in[45]
  PIN io_sram5_rw_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END io_sram5_rw_in[46]
  PIN io_sram5_rw_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 796.000 200.470 800.000 ;
    END
  END io_sram5_rw_in[47]
  PIN io_sram5_rw_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.840 500.000 177.440 ;
    END
  END io_sram5_rw_in[48]
  PIN io_sram5_rw_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END io_sram5_rw_in[49]
  PIN io_sram5_rw_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 796.000 248.770 800.000 ;
    END
  END io_sram5_rw_in[4]
  PIN io_sram5_rw_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_sram5_rw_in[50]
  PIN io_sram5_rw_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 360.440 500.000 361.040 ;
    END
  END io_sram5_rw_in[51]
  PIN io_sram5_rw_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END io_sram5_rw_in[52]
  PIN io_sram5_rw_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 796.000 458.070 800.000 ;
    END
  END io_sram5_rw_in[53]
  PIN io_sram5_rw_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 796.000 343.070 800.000 ;
    END
  END io_sram5_rw_in[54]
  PIN io_sram5_rw_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_sram5_rw_in[55]
  PIN io_sram5_rw_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END io_sram5_rw_in[56]
  PIN io_sram5_rw_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 796.000 67.070 800.000 ;
    END
  END io_sram5_rw_in[57]
  PIN io_sram5_rw_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END io_sram5_rw_in[58]
  PIN io_sram5_rw_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_sram5_rw_in[59]
  PIN io_sram5_rw_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_sram5_rw_in[5]
  PIN io_sram5_rw_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_sram5_rw_in[60]
  PIN io_sram5_rw_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 629.040 500.000 629.640 ;
    END
  END io_sram5_rw_in[61]
  PIN io_sram5_rw_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END io_sram5_rw_in[62]
  PIN io_sram5_rw_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_sram5_rw_in[63]
  PIN io_sram5_rw_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 136.040 500.000 136.640 ;
    END
  END io_sram5_rw_in[6]
  PIN io_sram5_rw_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END io_sram5_rw_in[7]
  PIN io_sram5_rw_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 23.840 500.000 24.440 ;
    END
  END io_sram5_rw_in[8]
  PIN io_sram5_rw_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 796.000 297.070 800.000 ;
    END
  END io_sram5_rw_in[9]
  PIN io_sram_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 516.840 500.000 517.440 ;
    END
  END io_sram_data[0]
  PIN io_sram_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 796.000 287.870 800.000 ;
    END
  END io_sram_data[10]
  PIN io_sram_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END io_sram_data[11]
  PIN io_sram_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 796.000 202.770 800.000 ;
    END
  END io_sram_data[12]
  PIN io_sram_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.040 500.000 442.640 ;
    END
  END io_sram_data[13]
  PIN io_sram_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 703.840 500.000 704.440 ;
    END
  END io_sram_data[14]
  PIN io_sram_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END io_sram_data[15]
  PIN io_sram_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END io_sram_data[16]
  PIN io_sram_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 796.000 50.970 800.000 ;
    END
  END io_sram_data[17]
  PIN io_sram_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END io_sram_data[18]
  PIN io_sram_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END io_sram_data[19]
  PIN io_sram_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 796.000 439.670 800.000 ;
    END
  END io_sram_data[1]
  PIN io_sram_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_sram_data[20]
  PIN io_sram_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 796.000 234.970 800.000 ;
    END
  END io_sram_data[21]
  PIN io_sram_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_sram_data[22]
  PIN io_sram_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 796.000 83.170 800.000 ;
    END
  END io_sram_data[23]
  PIN io_sram_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 496.440 500.000 497.040 ;
    END
  END io_sram_data[24]
  PIN io_sram_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 796.000 462.670 800.000 ;
    END
  END io_sram_data[25]
  PIN io_sram_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 796.000 23.370 800.000 ;
    END
  END io_sram_data[26]
  PIN io_sram_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 564.440 500.000 565.040 ;
    END
  END io_sram_data[27]
  PIN io_sram_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_sram_data[28]
  PIN io_sram_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END io_sram_data[29]
  PIN io_sram_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END io_sram_data[2]
  PIN io_sram_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 646.040 500.000 646.640 ;
    END
  END io_sram_data[30]
  PIN io_sram_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END io_sram_data[31]
  PIN io_sram_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 796.000 223.470 800.000 ;
    END
  END io_sram_data[32]
  PIN io_sram_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END io_sram_data[33]
  PIN io_sram_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END io_sram_data[34]
  PIN io_sram_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END io_sram_data[35]
  PIN io_sram_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END io_sram_data[36]
  PIN io_sram_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END io_sram_data[37]
  PIN io_sram_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 605.240 500.000 605.840 ;
    END
  END io_sram_data[38]
  PIN io_sram_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END io_sram_data[39]
  PIN io_sram_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 411.440 500.000 412.040 ;
    END
  END io_sram_data[3]
  PIN io_sram_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 258.440 500.000 259.040 ;
    END
  END io_sram_data[40]
  PIN io_sram_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END io_sram_data[41]
  PIN io_sram_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 581.440 500.000 582.040 ;
    END
  END io_sram_data[42]
  PIN io_sram_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END io_sram_data[43]
  PIN io_sram_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 796.000 179.770 800.000 ;
    END
  END io_sram_data[44]
  PIN io_sram_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END io_sram_data[45]
  PIN io_sram_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 796.000 354.570 800.000 ;
    END
  END io_sram_data[46]
  PIN io_sram_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END io_sram_data[47]
  PIN io_sram_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 707.240 500.000 707.840 ;
    END
  END io_sram_data[48]
  PIN io_sram_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END io_sram_data[49]
  PIN io_sram_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END io_sram_data[4]
  PIN io_sram_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_sram_data[50]
  PIN io_sram_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 724.240 500.000 724.840 ;
    END
  END io_sram_data[51]
  PIN io_sram_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END io_sram_data[52]
  PIN io_sram_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END io_sram_data[53]
  PIN io_sram_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END io_sram_data[54]
  PIN io_sram_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 537.240 500.000 537.840 ;
    END
  END io_sram_data[55]
  PIN io_sram_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END io_sram_data[56]
  PIN io_sram_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 255.040 500.000 255.640 ;
    END
  END io_sram_data[57]
  PIN io_sram_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END io_sram_data[58]
  PIN io_sram_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 796.000 269.470 800.000 ;
    END
  END io_sram_data[59]
  PIN io_sram_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END io_sram_data[5]
  PIN io_sram_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 796.000 168.270 800.000 ;
    END
  END io_sram_data[60]
  PIN io_sram_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END io_sram_data[61]
  PIN io_sram_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_sram_data[62]
  PIN io_sram_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END io_sram_data[63]
  PIN io_sram_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 796.000 428.170 800.000 ;
    END
  END io_sram_data[6]
  PIN io_sram_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 693.640 500.000 694.240 ;
    END
  END io_sram_data[7]
  PIN io_sram_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 796.000 163.670 800.000 ;
    END
  END io_sram_data[8]
  PIN io_sram_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_sram_data[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.040 500.000 408.640 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 788.800 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 788.800 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 788.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 788.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 788.800 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 788.800 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 788.885 ;
      LAYER met1 ;
        RECT 2.370 7.860 497.190 790.800 ;
      LAYER met2 ;
        RECT 2.400 795.720 4.410 796.125 ;
        RECT 5.250 795.720 6.710 796.125 ;
        RECT 7.550 795.720 9.010 796.125 ;
        RECT 9.850 795.720 11.310 796.125 ;
        RECT 12.150 795.720 13.610 796.125 ;
        RECT 14.450 795.720 15.910 796.125 ;
        RECT 16.750 795.720 18.210 796.125 ;
        RECT 19.050 795.720 20.510 796.125 ;
        RECT 21.350 795.720 22.810 796.125 ;
        RECT 23.650 795.720 25.110 796.125 ;
        RECT 25.950 795.720 27.410 796.125 ;
        RECT 28.250 795.720 29.710 796.125 ;
        RECT 30.550 795.720 34.310 796.125 ;
        RECT 35.150 795.720 36.610 796.125 ;
        RECT 37.450 795.720 38.910 796.125 ;
        RECT 39.750 795.720 41.210 796.125 ;
        RECT 42.050 795.720 43.510 796.125 ;
        RECT 44.350 795.720 45.810 796.125 ;
        RECT 46.650 795.720 48.110 796.125 ;
        RECT 48.950 795.720 50.410 796.125 ;
        RECT 51.250 795.720 52.710 796.125 ;
        RECT 53.550 795.720 55.010 796.125 ;
        RECT 55.850 795.720 57.310 796.125 ;
        RECT 58.150 795.720 59.610 796.125 ;
        RECT 60.450 795.720 64.210 796.125 ;
        RECT 65.050 795.720 66.510 796.125 ;
        RECT 67.350 795.720 68.810 796.125 ;
        RECT 69.650 795.720 71.110 796.125 ;
        RECT 71.950 795.720 73.410 796.125 ;
        RECT 74.250 795.720 75.710 796.125 ;
        RECT 76.550 795.720 78.010 796.125 ;
        RECT 78.850 795.720 80.310 796.125 ;
        RECT 81.150 795.720 82.610 796.125 ;
        RECT 83.450 795.720 84.910 796.125 ;
        RECT 85.750 795.720 87.210 796.125 ;
        RECT 88.050 795.720 89.510 796.125 ;
        RECT 90.350 795.720 94.110 796.125 ;
        RECT 94.950 795.720 96.410 796.125 ;
        RECT 97.250 795.720 98.710 796.125 ;
        RECT 99.550 795.720 101.010 796.125 ;
        RECT 101.850 795.720 103.310 796.125 ;
        RECT 104.150 795.720 105.610 796.125 ;
        RECT 106.450 795.720 107.910 796.125 ;
        RECT 108.750 795.720 110.210 796.125 ;
        RECT 111.050 795.720 112.510 796.125 ;
        RECT 113.350 795.720 114.810 796.125 ;
        RECT 115.650 795.720 117.110 796.125 ;
        RECT 117.950 795.720 119.410 796.125 ;
        RECT 120.250 795.720 124.010 796.125 ;
        RECT 124.850 795.720 126.310 796.125 ;
        RECT 127.150 795.720 128.610 796.125 ;
        RECT 129.450 795.720 130.910 796.125 ;
        RECT 131.750 795.720 133.210 796.125 ;
        RECT 134.050 795.720 135.510 796.125 ;
        RECT 136.350 795.720 137.810 796.125 ;
        RECT 138.650 795.720 140.110 796.125 ;
        RECT 140.950 795.720 142.410 796.125 ;
        RECT 143.250 795.720 144.710 796.125 ;
        RECT 145.550 795.720 147.010 796.125 ;
        RECT 147.850 795.720 149.310 796.125 ;
        RECT 150.150 795.720 151.610 796.125 ;
        RECT 152.450 795.720 156.210 796.125 ;
        RECT 157.050 795.720 158.510 796.125 ;
        RECT 159.350 795.720 160.810 796.125 ;
        RECT 161.650 795.720 163.110 796.125 ;
        RECT 163.950 795.720 165.410 796.125 ;
        RECT 166.250 795.720 167.710 796.125 ;
        RECT 168.550 795.720 170.010 796.125 ;
        RECT 170.850 795.720 172.310 796.125 ;
        RECT 173.150 795.720 174.610 796.125 ;
        RECT 175.450 795.720 176.910 796.125 ;
        RECT 177.750 795.720 179.210 796.125 ;
        RECT 180.050 795.720 181.510 796.125 ;
        RECT 182.350 795.720 186.110 796.125 ;
        RECT 186.950 795.720 188.410 796.125 ;
        RECT 189.250 795.720 190.710 796.125 ;
        RECT 191.550 795.720 193.010 796.125 ;
        RECT 193.850 795.720 195.310 796.125 ;
        RECT 196.150 795.720 197.610 796.125 ;
        RECT 198.450 795.720 199.910 796.125 ;
        RECT 200.750 795.720 202.210 796.125 ;
        RECT 203.050 795.720 204.510 796.125 ;
        RECT 205.350 795.720 206.810 796.125 ;
        RECT 207.650 795.720 209.110 796.125 ;
        RECT 209.950 795.720 211.410 796.125 ;
        RECT 212.250 795.720 216.010 796.125 ;
        RECT 216.850 795.720 218.310 796.125 ;
        RECT 219.150 795.720 220.610 796.125 ;
        RECT 221.450 795.720 222.910 796.125 ;
        RECT 223.750 795.720 225.210 796.125 ;
        RECT 226.050 795.720 227.510 796.125 ;
        RECT 228.350 795.720 229.810 796.125 ;
        RECT 230.650 795.720 232.110 796.125 ;
        RECT 232.950 795.720 234.410 796.125 ;
        RECT 235.250 795.720 236.710 796.125 ;
        RECT 237.550 795.720 239.010 796.125 ;
        RECT 239.850 795.720 241.310 796.125 ;
        RECT 242.150 795.720 245.910 796.125 ;
        RECT 246.750 795.720 248.210 796.125 ;
        RECT 249.050 795.720 250.510 796.125 ;
        RECT 251.350 795.720 252.810 796.125 ;
        RECT 253.650 795.720 255.110 796.125 ;
        RECT 255.950 795.720 257.410 796.125 ;
        RECT 258.250 795.720 259.710 796.125 ;
        RECT 260.550 795.720 262.010 796.125 ;
        RECT 262.850 795.720 264.310 796.125 ;
        RECT 265.150 795.720 266.610 796.125 ;
        RECT 267.450 795.720 268.910 796.125 ;
        RECT 269.750 795.720 271.210 796.125 ;
        RECT 272.050 795.720 275.810 796.125 ;
        RECT 276.650 795.720 278.110 796.125 ;
        RECT 278.950 795.720 280.410 796.125 ;
        RECT 281.250 795.720 282.710 796.125 ;
        RECT 283.550 795.720 285.010 796.125 ;
        RECT 285.850 795.720 287.310 796.125 ;
        RECT 288.150 795.720 289.610 796.125 ;
        RECT 290.450 795.720 291.910 796.125 ;
        RECT 292.750 795.720 294.210 796.125 ;
        RECT 295.050 795.720 296.510 796.125 ;
        RECT 297.350 795.720 298.810 796.125 ;
        RECT 299.650 795.720 301.110 796.125 ;
        RECT 301.950 795.720 305.710 796.125 ;
        RECT 306.550 795.720 308.010 796.125 ;
        RECT 308.850 795.720 310.310 796.125 ;
        RECT 311.150 795.720 312.610 796.125 ;
        RECT 313.450 795.720 314.910 796.125 ;
        RECT 315.750 795.720 317.210 796.125 ;
        RECT 318.050 795.720 319.510 796.125 ;
        RECT 320.350 795.720 321.810 796.125 ;
        RECT 322.650 795.720 324.110 796.125 ;
        RECT 324.950 795.720 326.410 796.125 ;
        RECT 327.250 795.720 328.710 796.125 ;
        RECT 329.550 795.720 331.010 796.125 ;
        RECT 331.850 795.720 335.610 796.125 ;
        RECT 336.450 795.720 337.910 796.125 ;
        RECT 338.750 795.720 340.210 796.125 ;
        RECT 341.050 795.720 342.510 796.125 ;
        RECT 343.350 795.720 344.810 796.125 ;
        RECT 345.650 795.720 347.110 796.125 ;
        RECT 347.950 795.720 349.410 796.125 ;
        RECT 350.250 795.720 351.710 796.125 ;
        RECT 352.550 795.720 354.010 796.125 ;
        RECT 354.850 795.720 356.310 796.125 ;
        RECT 357.150 795.720 358.610 796.125 ;
        RECT 359.450 795.720 360.910 796.125 ;
        RECT 361.750 795.720 365.510 796.125 ;
        RECT 366.350 795.720 367.810 796.125 ;
        RECT 368.650 795.720 370.110 796.125 ;
        RECT 370.950 795.720 372.410 796.125 ;
        RECT 373.250 795.720 374.710 796.125 ;
        RECT 375.550 795.720 377.010 796.125 ;
        RECT 377.850 795.720 379.310 796.125 ;
        RECT 380.150 795.720 381.610 796.125 ;
        RECT 382.450 795.720 383.910 796.125 ;
        RECT 384.750 795.720 386.210 796.125 ;
        RECT 387.050 795.720 388.510 796.125 ;
        RECT 389.350 795.720 390.810 796.125 ;
        RECT 391.650 795.720 395.410 796.125 ;
        RECT 396.250 795.720 397.710 796.125 ;
        RECT 398.550 795.720 400.010 796.125 ;
        RECT 400.850 795.720 402.310 796.125 ;
        RECT 403.150 795.720 404.610 796.125 ;
        RECT 405.450 795.720 406.910 796.125 ;
        RECT 407.750 795.720 409.210 796.125 ;
        RECT 410.050 795.720 411.510 796.125 ;
        RECT 412.350 795.720 413.810 796.125 ;
        RECT 414.650 795.720 416.110 796.125 ;
        RECT 416.950 795.720 418.410 796.125 ;
        RECT 419.250 795.720 420.710 796.125 ;
        RECT 421.550 795.720 425.310 796.125 ;
        RECT 426.150 795.720 427.610 796.125 ;
        RECT 428.450 795.720 429.910 796.125 ;
        RECT 430.750 795.720 432.210 796.125 ;
        RECT 433.050 795.720 434.510 796.125 ;
        RECT 435.350 795.720 436.810 796.125 ;
        RECT 437.650 795.720 439.110 796.125 ;
        RECT 439.950 795.720 441.410 796.125 ;
        RECT 442.250 795.720 443.710 796.125 ;
        RECT 444.550 795.720 446.010 796.125 ;
        RECT 446.850 795.720 448.310 796.125 ;
        RECT 449.150 795.720 450.610 796.125 ;
        RECT 451.450 795.720 455.210 796.125 ;
        RECT 456.050 795.720 457.510 796.125 ;
        RECT 458.350 795.720 459.810 796.125 ;
        RECT 460.650 795.720 462.110 796.125 ;
        RECT 462.950 795.720 464.410 796.125 ;
        RECT 465.250 795.720 466.710 796.125 ;
        RECT 467.550 795.720 469.010 796.125 ;
        RECT 469.850 795.720 471.310 796.125 ;
        RECT 472.150 795.720 473.610 796.125 ;
        RECT 474.450 795.720 475.910 796.125 ;
        RECT 476.750 795.720 478.210 796.125 ;
        RECT 479.050 795.720 480.510 796.125 ;
        RECT 481.350 795.720 485.110 796.125 ;
        RECT 485.950 795.720 487.410 796.125 ;
        RECT 488.250 795.720 489.710 796.125 ;
        RECT 490.550 795.720 492.010 796.125 ;
        RECT 492.850 795.720 494.310 796.125 ;
        RECT 495.150 795.720 496.610 796.125 ;
        RECT 2.400 4.280 497.160 795.720 ;
        RECT 2.950 3.555 4.410 4.280 ;
        RECT 5.250 3.555 6.710 4.280 ;
        RECT 7.550 3.555 9.010 4.280 ;
        RECT 9.850 3.555 11.310 4.280 ;
        RECT 12.150 3.555 13.610 4.280 ;
        RECT 14.450 3.555 15.910 4.280 ;
        RECT 16.750 3.555 18.210 4.280 ;
        RECT 19.050 3.555 20.510 4.280 ;
        RECT 21.350 3.555 22.810 4.280 ;
        RECT 23.650 3.555 25.110 4.280 ;
        RECT 25.950 3.555 27.410 4.280 ;
        RECT 28.250 3.555 29.710 4.280 ;
        RECT 30.550 3.555 34.310 4.280 ;
        RECT 35.150 3.555 36.610 4.280 ;
        RECT 37.450 3.555 38.910 4.280 ;
        RECT 39.750 3.555 41.210 4.280 ;
        RECT 42.050 3.555 43.510 4.280 ;
        RECT 44.350 3.555 45.810 4.280 ;
        RECT 46.650 3.555 48.110 4.280 ;
        RECT 48.950 3.555 50.410 4.280 ;
        RECT 51.250 3.555 52.710 4.280 ;
        RECT 53.550 3.555 55.010 4.280 ;
        RECT 55.850 3.555 57.310 4.280 ;
        RECT 58.150 3.555 59.610 4.280 ;
        RECT 60.450 3.555 64.210 4.280 ;
        RECT 65.050 3.555 66.510 4.280 ;
        RECT 67.350 3.555 68.810 4.280 ;
        RECT 69.650 3.555 71.110 4.280 ;
        RECT 71.950 3.555 73.410 4.280 ;
        RECT 74.250 3.555 75.710 4.280 ;
        RECT 76.550 3.555 78.010 4.280 ;
        RECT 78.850 3.555 80.310 4.280 ;
        RECT 81.150 3.555 82.610 4.280 ;
        RECT 83.450 3.555 84.910 4.280 ;
        RECT 85.750 3.555 87.210 4.280 ;
        RECT 88.050 3.555 89.510 4.280 ;
        RECT 90.350 3.555 94.110 4.280 ;
        RECT 94.950 3.555 96.410 4.280 ;
        RECT 97.250 3.555 98.710 4.280 ;
        RECT 99.550 3.555 101.010 4.280 ;
        RECT 101.850 3.555 103.310 4.280 ;
        RECT 104.150 3.555 105.610 4.280 ;
        RECT 106.450 3.555 107.910 4.280 ;
        RECT 108.750 3.555 110.210 4.280 ;
        RECT 111.050 3.555 112.510 4.280 ;
        RECT 113.350 3.555 114.810 4.280 ;
        RECT 115.650 3.555 117.110 4.280 ;
        RECT 117.950 3.555 119.410 4.280 ;
        RECT 120.250 3.555 124.010 4.280 ;
        RECT 124.850 3.555 126.310 4.280 ;
        RECT 127.150 3.555 128.610 4.280 ;
        RECT 129.450 3.555 130.910 4.280 ;
        RECT 131.750 3.555 133.210 4.280 ;
        RECT 134.050 3.555 135.510 4.280 ;
        RECT 136.350 3.555 137.810 4.280 ;
        RECT 138.650 3.555 140.110 4.280 ;
        RECT 140.950 3.555 142.410 4.280 ;
        RECT 143.250 3.555 144.710 4.280 ;
        RECT 145.550 3.555 147.010 4.280 ;
        RECT 147.850 3.555 149.310 4.280 ;
        RECT 150.150 3.555 153.910 4.280 ;
        RECT 154.750 3.555 156.210 4.280 ;
        RECT 157.050 3.555 158.510 4.280 ;
        RECT 159.350 3.555 160.810 4.280 ;
        RECT 161.650 3.555 163.110 4.280 ;
        RECT 163.950 3.555 165.410 4.280 ;
        RECT 166.250 3.555 167.710 4.280 ;
        RECT 168.550 3.555 170.010 4.280 ;
        RECT 170.850 3.555 172.310 4.280 ;
        RECT 173.150 3.555 174.610 4.280 ;
        RECT 175.450 3.555 176.910 4.280 ;
        RECT 177.750 3.555 179.210 4.280 ;
        RECT 180.050 3.555 183.810 4.280 ;
        RECT 184.650 3.555 186.110 4.280 ;
        RECT 186.950 3.555 188.410 4.280 ;
        RECT 189.250 3.555 190.710 4.280 ;
        RECT 191.550 3.555 193.010 4.280 ;
        RECT 193.850 3.555 195.310 4.280 ;
        RECT 196.150 3.555 197.610 4.280 ;
        RECT 198.450 3.555 199.910 4.280 ;
        RECT 200.750 3.555 202.210 4.280 ;
        RECT 203.050 3.555 204.510 4.280 ;
        RECT 205.350 3.555 206.810 4.280 ;
        RECT 207.650 3.555 209.110 4.280 ;
        RECT 209.950 3.555 213.710 4.280 ;
        RECT 214.550 3.555 216.010 4.280 ;
        RECT 216.850 3.555 218.310 4.280 ;
        RECT 219.150 3.555 220.610 4.280 ;
        RECT 221.450 3.555 222.910 4.280 ;
        RECT 223.750 3.555 225.210 4.280 ;
        RECT 226.050 3.555 227.510 4.280 ;
        RECT 228.350 3.555 229.810 4.280 ;
        RECT 230.650 3.555 232.110 4.280 ;
        RECT 232.950 3.555 234.410 4.280 ;
        RECT 235.250 3.555 236.710 4.280 ;
        RECT 237.550 3.555 239.010 4.280 ;
        RECT 239.850 3.555 243.610 4.280 ;
        RECT 244.450 3.555 245.910 4.280 ;
        RECT 246.750 3.555 248.210 4.280 ;
        RECT 249.050 3.555 250.510 4.280 ;
        RECT 251.350 3.555 252.810 4.280 ;
        RECT 253.650 3.555 255.110 4.280 ;
        RECT 255.950 3.555 257.410 4.280 ;
        RECT 258.250 3.555 259.710 4.280 ;
        RECT 260.550 3.555 262.010 4.280 ;
        RECT 262.850 3.555 264.310 4.280 ;
        RECT 265.150 3.555 266.610 4.280 ;
        RECT 267.450 3.555 268.910 4.280 ;
        RECT 269.750 3.555 273.510 4.280 ;
        RECT 274.350 3.555 275.810 4.280 ;
        RECT 276.650 3.555 278.110 4.280 ;
        RECT 278.950 3.555 280.410 4.280 ;
        RECT 281.250 3.555 282.710 4.280 ;
        RECT 283.550 3.555 285.010 4.280 ;
        RECT 285.850 3.555 287.310 4.280 ;
        RECT 288.150 3.555 289.610 4.280 ;
        RECT 290.450 3.555 291.910 4.280 ;
        RECT 292.750 3.555 294.210 4.280 ;
        RECT 295.050 3.555 296.510 4.280 ;
        RECT 297.350 3.555 298.810 4.280 ;
        RECT 299.650 3.555 303.410 4.280 ;
        RECT 304.250 3.555 305.710 4.280 ;
        RECT 306.550 3.555 308.010 4.280 ;
        RECT 308.850 3.555 310.310 4.280 ;
        RECT 311.150 3.555 312.610 4.280 ;
        RECT 313.450 3.555 314.910 4.280 ;
        RECT 315.750 3.555 317.210 4.280 ;
        RECT 318.050 3.555 319.510 4.280 ;
        RECT 320.350 3.555 321.810 4.280 ;
        RECT 322.650 3.555 324.110 4.280 ;
        RECT 324.950 3.555 326.410 4.280 ;
        RECT 327.250 3.555 328.710 4.280 ;
        RECT 329.550 3.555 333.310 4.280 ;
        RECT 334.150 3.555 335.610 4.280 ;
        RECT 336.450 3.555 337.910 4.280 ;
        RECT 338.750 3.555 340.210 4.280 ;
        RECT 341.050 3.555 342.510 4.280 ;
        RECT 343.350 3.555 344.810 4.280 ;
        RECT 345.650 3.555 347.110 4.280 ;
        RECT 347.950 3.555 349.410 4.280 ;
        RECT 350.250 3.555 351.710 4.280 ;
        RECT 352.550 3.555 354.010 4.280 ;
        RECT 354.850 3.555 356.310 4.280 ;
        RECT 357.150 3.555 358.610 4.280 ;
        RECT 359.450 3.555 363.210 4.280 ;
        RECT 364.050 3.555 365.510 4.280 ;
        RECT 366.350 3.555 367.810 4.280 ;
        RECT 368.650 3.555 370.110 4.280 ;
        RECT 370.950 3.555 372.410 4.280 ;
        RECT 373.250 3.555 374.710 4.280 ;
        RECT 375.550 3.555 377.010 4.280 ;
        RECT 377.850 3.555 379.310 4.280 ;
        RECT 380.150 3.555 381.610 4.280 ;
        RECT 382.450 3.555 383.910 4.280 ;
        RECT 384.750 3.555 386.210 4.280 ;
        RECT 387.050 3.555 388.510 4.280 ;
        RECT 389.350 3.555 393.110 4.280 ;
        RECT 393.950 3.555 395.410 4.280 ;
        RECT 396.250 3.555 397.710 4.280 ;
        RECT 398.550 3.555 400.010 4.280 ;
        RECT 400.850 3.555 402.310 4.280 ;
        RECT 403.150 3.555 404.610 4.280 ;
        RECT 405.450 3.555 406.910 4.280 ;
        RECT 407.750 3.555 409.210 4.280 ;
        RECT 410.050 3.555 411.510 4.280 ;
        RECT 412.350 3.555 413.810 4.280 ;
        RECT 414.650 3.555 416.110 4.280 ;
        RECT 416.950 3.555 418.410 4.280 ;
        RECT 419.250 3.555 423.010 4.280 ;
        RECT 423.850 3.555 425.310 4.280 ;
        RECT 426.150 3.555 427.610 4.280 ;
        RECT 428.450 3.555 429.910 4.280 ;
        RECT 430.750 3.555 432.210 4.280 ;
        RECT 433.050 3.555 434.510 4.280 ;
        RECT 435.350 3.555 436.810 4.280 ;
        RECT 437.650 3.555 439.110 4.280 ;
        RECT 439.950 3.555 441.410 4.280 ;
        RECT 442.250 3.555 443.710 4.280 ;
        RECT 444.550 3.555 446.010 4.280 ;
        RECT 446.850 3.555 448.310 4.280 ;
        RECT 449.150 3.555 452.910 4.280 ;
        RECT 453.750 3.555 455.210 4.280 ;
        RECT 456.050 3.555 457.510 4.280 ;
        RECT 458.350 3.555 459.810 4.280 ;
        RECT 460.650 3.555 462.110 4.280 ;
        RECT 462.950 3.555 464.410 4.280 ;
        RECT 465.250 3.555 466.710 4.280 ;
        RECT 467.550 3.555 469.010 4.280 ;
        RECT 469.850 3.555 471.310 4.280 ;
        RECT 472.150 3.555 473.610 4.280 ;
        RECT 474.450 3.555 475.910 4.280 ;
        RECT 476.750 3.555 478.210 4.280 ;
        RECT 479.050 3.555 482.810 4.280 ;
        RECT 483.650 3.555 485.110 4.280 ;
        RECT 485.950 3.555 487.410 4.280 ;
        RECT 488.250 3.555 489.710 4.280 ;
        RECT 490.550 3.555 492.010 4.280 ;
        RECT 492.850 3.555 494.310 4.280 ;
        RECT 495.150 3.555 496.610 4.280 ;
      LAYER met3 ;
        RECT 4.400 795.240 495.600 796.105 ;
        RECT 4.000 793.240 496.000 795.240 ;
        RECT 4.400 791.840 495.600 793.240 ;
        RECT 4.000 789.840 496.000 791.840 ;
        RECT 4.400 788.440 495.600 789.840 ;
        RECT 4.000 786.440 496.000 788.440 ;
        RECT 4.400 785.040 495.600 786.440 ;
        RECT 4.000 783.040 496.000 785.040 ;
        RECT 4.400 781.640 495.600 783.040 ;
        RECT 4.000 779.640 496.000 781.640 ;
        RECT 4.400 778.240 495.600 779.640 ;
        RECT 4.000 776.240 496.000 778.240 ;
        RECT 4.400 774.840 496.000 776.240 ;
        RECT 4.000 772.840 496.000 774.840 ;
        RECT 4.400 771.440 495.600 772.840 ;
        RECT 4.000 769.440 496.000 771.440 ;
        RECT 4.400 768.040 495.600 769.440 ;
        RECT 4.000 766.040 496.000 768.040 ;
        RECT 4.400 764.640 495.600 766.040 ;
        RECT 4.000 762.640 496.000 764.640 ;
        RECT 4.400 761.240 495.600 762.640 ;
        RECT 4.000 759.240 496.000 761.240 ;
        RECT 4.400 757.840 495.600 759.240 ;
        RECT 4.000 755.840 496.000 757.840 ;
        RECT 4.000 754.440 495.600 755.840 ;
        RECT 4.000 752.440 496.000 754.440 ;
        RECT 4.400 751.040 495.600 752.440 ;
        RECT 4.000 749.040 496.000 751.040 ;
        RECT 4.400 747.640 495.600 749.040 ;
        RECT 4.000 745.640 496.000 747.640 ;
        RECT 4.400 744.240 495.600 745.640 ;
        RECT 4.000 742.240 496.000 744.240 ;
        RECT 4.400 740.840 495.600 742.240 ;
        RECT 4.000 738.840 496.000 740.840 ;
        RECT 4.400 737.440 495.600 738.840 ;
        RECT 4.000 735.440 496.000 737.440 ;
        RECT 4.400 734.040 495.600 735.440 ;
        RECT 4.000 732.040 496.000 734.040 ;
        RECT 4.400 730.640 496.000 732.040 ;
        RECT 4.000 728.640 496.000 730.640 ;
        RECT 4.400 727.240 495.600 728.640 ;
        RECT 4.000 725.240 496.000 727.240 ;
        RECT 4.400 723.840 495.600 725.240 ;
        RECT 4.000 721.840 496.000 723.840 ;
        RECT 4.400 720.440 495.600 721.840 ;
        RECT 4.000 718.440 496.000 720.440 ;
        RECT 4.400 717.040 495.600 718.440 ;
        RECT 4.000 715.040 496.000 717.040 ;
        RECT 4.400 713.640 495.600 715.040 ;
        RECT 4.000 711.640 496.000 713.640 ;
        RECT 4.000 710.240 495.600 711.640 ;
        RECT 4.000 708.240 496.000 710.240 ;
        RECT 4.400 706.840 495.600 708.240 ;
        RECT 4.000 704.840 496.000 706.840 ;
        RECT 4.400 703.440 495.600 704.840 ;
        RECT 4.000 701.440 496.000 703.440 ;
        RECT 4.400 700.040 495.600 701.440 ;
        RECT 4.000 698.040 496.000 700.040 ;
        RECT 4.400 696.640 495.600 698.040 ;
        RECT 4.000 694.640 496.000 696.640 ;
        RECT 4.400 693.240 495.600 694.640 ;
        RECT 4.000 691.240 496.000 693.240 ;
        RECT 4.400 689.840 495.600 691.240 ;
        RECT 4.000 687.840 496.000 689.840 ;
        RECT 4.400 686.440 496.000 687.840 ;
        RECT 4.000 684.440 496.000 686.440 ;
        RECT 4.400 683.040 495.600 684.440 ;
        RECT 4.000 681.040 496.000 683.040 ;
        RECT 4.400 679.640 495.600 681.040 ;
        RECT 4.000 677.640 496.000 679.640 ;
        RECT 4.400 676.240 495.600 677.640 ;
        RECT 4.000 674.240 496.000 676.240 ;
        RECT 4.400 672.840 495.600 674.240 ;
        RECT 4.000 670.840 496.000 672.840 ;
        RECT 4.400 669.440 495.600 670.840 ;
        RECT 4.000 667.440 496.000 669.440 ;
        RECT 4.000 666.040 495.600 667.440 ;
        RECT 4.000 664.040 496.000 666.040 ;
        RECT 4.400 662.640 495.600 664.040 ;
        RECT 4.000 660.640 496.000 662.640 ;
        RECT 4.400 659.240 495.600 660.640 ;
        RECT 4.000 657.240 496.000 659.240 ;
        RECT 4.400 655.840 495.600 657.240 ;
        RECT 4.000 653.840 496.000 655.840 ;
        RECT 4.400 652.440 495.600 653.840 ;
        RECT 4.000 650.440 496.000 652.440 ;
        RECT 4.400 649.040 495.600 650.440 ;
        RECT 4.000 647.040 496.000 649.040 ;
        RECT 4.400 645.640 495.600 647.040 ;
        RECT 4.000 643.640 496.000 645.640 ;
        RECT 4.400 642.240 496.000 643.640 ;
        RECT 4.000 640.240 496.000 642.240 ;
        RECT 4.400 638.840 495.600 640.240 ;
        RECT 4.000 636.840 496.000 638.840 ;
        RECT 4.400 635.440 495.600 636.840 ;
        RECT 4.000 633.440 496.000 635.440 ;
        RECT 4.400 632.040 495.600 633.440 ;
        RECT 4.000 630.040 496.000 632.040 ;
        RECT 4.400 628.640 495.600 630.040 ;
        RECT 4.000 626.640 496.000 628.640 ;
        RECT 4.400 625.240 495.600 626.640 ;
        RECT 4.000 623.240 496.000 625.240 ;
        RECT 4.000 621.840 495.600 623.240 ;
        RECT 4.000 619.840 496.000 621.840 ;
        RECT 4.400 618.440 495.600 619.840 ;
        RECT 4.000 616.440 496.000 618.440 ;
        RECT 4.400 615.040 495.600 616.440 ;
        RECT 4.000 613.040 496.000 615.040 ;
        RECT 4.400 611.640 495.600 613.040 ;
        RECT 4.000 609.640 496.000 611.640 ;
        RECT 4.400 608.240 495.600 609.640 ;
        RECT 4.000 606.240 496.000 608.240 ;
        RECT 4.400 604.840 495.600 606.240 ;
        RECT 4.000 602.840 496.000 604.840 ;
        RECT 4.400 601.440 495.600 602.840 ;
        RECT 4.000 599.440 496.000 601.440 ;
        RECT 4.400 598.040 496.000 599.440 ;
        RECT 4.000 596.040 496.000 598.040 ;
        RECT 4.400 594.640 495.600 596.040 ;
        RECT 4.000 592.640 496.000 594.640 ;
        RECT 4.400 591.240 495.600 592.640 ;
        RECT 4.000 589.240 496.000 591.240 ;
        RECT 4.400 587.840 495.600 589.240 ;
        RECT 4.000 585.840 496.000 587.840 ;
        RECT 4.400 584.440 495.600 585.840 ;
        RECT 4.000 582.440 496.000 584.440 ;
        RECT 4.400 581.040 495.600 582.440 ;
        RECT 4.000 579.040 496.000 581.040 ;
        RECT 4.000 577.640 495.600 579.040 ;
        RECT 4.000 575.640 496.000 577.640 ;
        RECT 4.400 574.240 495.600 575.640 ;
        RECT 4.000 572.240 496.000 574.240 ;
        RECT 4.400 570.840 495.600 572.240 ;
        RECT 4.000 568.840 496.000 570.840 ;
        RECT 4.400 567.440 495.600 568.840 ;
        RECT 4.000 565.440 496.000 567.440 ;
        RECT 4.400 564.040 495.600 565.440 ;
        RECT 4.000 562.040 496.000 564.040 ;
        RECT 4.400 560.640 495.600 562.040 ;
        RECT 4.000 558.640 496.000 560.640 ;
        RECT 4.400 557.240 495.600 558.640 ;
        RECT 4.000 555.240 496.000 557.240 ;
        RECT 4.400 553.840 496.000 555.240 ;
        RECT 4.000 551.840 496.000 553.840 ;
        RECT 4.400 550.440 495.600 551.840 ;
        RECT 4.000 548.440 496.000 550.440 ;
        RECT 4.400 547.040 495.600 548.440 ;
        RECT 4.000 545.040 496.000 547.040 ;
        RECT 4.400 543.640 495.600 545.040 ;
        RECT 4.000 541.640 496.000 543.640 ;
        RECT 4.400 540.240 495.600 541.640 ;
        RECT 4.000 538.240 496.000 540.240 ;
        RECT 4.400 536.840 495.600 538.240 ;
        RECT 4.000 534.840 496.000 536.840 ;
        RECT 4.000 533.440 495.600 534.840 ;
        RECT 4.000 531.440 496.000 533.440 ;
        RECT 4.400 530.040 495.600 531.440 ;
        RECT 4.000 528.040 496.000 530.040 ;
        RECT 4.400 526.640 495.600 528.040 ;
        RECT 4.000 524.640 496.000 526.640 ;
        RECT 4.400 523.240 495.600 524.640 ;
        RECT 4.000 521.240 496.000 523.240 ;
        RECT 4.400 519.840 495.600 521.240 ;
        RECT 4.000 517.840 496.000 519.840 ;
        RECT 4.400 516.440 495.600 517.840 ;
        RECT 4.000 514.440 496.000 516.440 ;
        RECT 4.400 513.040 495.600 514.440 ;
        RECT 4.000 511.040 496.000 513.040 ;
        RECT 4.400 509.640 496.000 511.040 ;
        RECT 4.000 507.640 496.000 509.640 ;
        RECT 4.400 506.240 495.600 507.640 ;
        RECT 4.000 504.240 496.000 506.240 ;
        RECT 4.400 502.840 495.600 504.240 ;
        RECT 4.000 500.840 496.000 502.840 ;
        RECT 4.400 499.440 495.600 500.840 ;
        RECT 4.000 497.440 496.000 499.440 ;
        RECT 4.400 496.040 495.600 497.440 ;
        RECT 4.000 494.040 496.000 496.040 ;
        RECT 4.400 492.640 495.600 494.040 ;
        RECT 4.000 490.640 496.000 492.640 ;
        RECT 4.000 489.240 495.600 490.640 ;
        RECT 4.000 487.240 496.000 489.240 ;
        RECT 4.400 485.840 495.600 487.240 ;
        RECT 4.000 483.840 496.000 485.840 ;
        RECT 4.400 482.440 495.600 483.840 ;
        RECT 4.000 480.440 496.000 482.440 ;
        RECT 4.400 479.040 495.600 480.440 ;
        RECT 4.000 477.040 496.000 479.040 ;
        RECT 4.400 475.640 495.600 477.040 ;
        RECT 4.000 473.640 496.000 475.640 ;
        RECT 4.400 472.240 495.600 473.640 ;
        RECT 4.000 470.240 496.000 472.240 ;
        RECT 4.400 468.840 495.600 470.240 ;
        RECT 4.000 466.840 496.000 468.840 ;
        RECT 4.400 465.440 496.000 466.840 ;
        RECT 4.000 463.440 496.000 465.440 ;
        RECT 4.400 462.040 495.600 463.440 ;
        RECT 4.000 460.040 496.000 462.040 ;
        RECT 4.400 458.640 495.600 460.040 ;
        RECT 4.000 456.640 496.000 458.640 ;
        RECT 4.400 455.240 495.600 456.640 ;
        RECT 4.000 453.240 496.000 455.240 ;
        RECT 4.400 451.840 495.600 453.240 ;
        RECT 4.000 449.840 496.000 451.840 ;
        RECT 4.400 448.440 495.600 449.840 ;
        RECT 4.000 446.440 496.000 448.440 ;
        RECT 4.000 445.040 495.600 446.440 ;
        RECT 4.000 443.040 496.000 445.040 ;
        RECT 4.400 441.640 495.600 443.040 ;
        RECT 4.000 439.640 496.000 441.640 ;
        RECT 4.400 438.240 495.600 439.640 ;
        RECT 4.000 436.240 496.000 438.240 ;
        RECT 4.400 434.840 495.600 436.240 ;
        RECT 4.000 432.840 496.000 434.840 ;
        RECT 4.400 431.440 495.600 432.840 ;
        RECT 4.000 429.440 496.000 431.440 ;
        RECT 4.400 428.040 495.600 429.440 ;
        RECT 4.000 426.040 496.000 428.040 ;
        RECT 4.400 424.640 495.600 426.040 ;
        RECT 4.000 422.640 496.000 424.640 ;
        RECT 4.400 421.240 496.000 422.640 ;
        RECT 4.000 419.240 496.000 421.240 ;
        RECT 4.400 417.840 495.600 419.240 ;
        RECT 4.000 415.840 496.000 417.840 ;
        RECT 4.400 414.440 495.600 415.840 ;
        RECT 4.000 412.440 496.000 414.440 ;
        RECT 4.400 411.040 495.600 412.440 ;
        RECT 4.000 409.040 496.000 411.040 ;
        RECT 4.400 407.640 495.600 409.040 ;
        RECT 4.000 405.640 496.000 407.640 ;
        RECT 4.400 404.240 495.600 405.640 ;
        RECT 4.000 402.240 496.000 404.240 ;
        RECT 4.000 400.840 495.600 402.240 ;
        RECT 4.000 398.840 496.000 400.840 ;
        RECT 4.400 397.440 495.600 398.840 ;
        RECT 4.000 395.440 496.000 397.440 ;
        RECT 4.400 394.040 495.600 395.440 ;
        RECT 4.000 392.040 496.000 394.040 ;
        RECT 4.400 390.640 495.600 392.040 ;
        RECT 4.000 388.640 496.000 390.640 ;
        RECT 4.400 387.240 495.600 388.640 ;
        RECT 4.000 385.240 496.000 387.240 ;
        RECT 4.400 383.840 495.600 385.240 ;
        RECT 4.000 381.840 496.000 383.840 ;
        RECT 4.400 380.440 495.600 381.840 ;
        RECT 4.000 378.440 496.000 380.440 ;
        RECT 4.400 377.040 496.000 378.440 ;
        RECT 4.000 375.040 496.000 377.040 ;
        RECT 4.400 373.640 495.600 375.040 ;
        RECT 4.000 371.640 496.000 373.640 ;
        RECT 4.400 370.240 495.600 371.640 ;
        RECT 4.000 368.240 496.000 370.240 ;
        RECT 4.400 366.840 495.600 368.240 ;
        RECT 4.000 364.840 496.000 366.840 ;
        RECT 4.400 363.440 495.600 364.840 ;
        RECT 4.000 361.440 496.000 363.440 ;
        RECT 4.400 360.040 495.600 361.440 ;
        RECT 4.000 358.040 496.000 360.040 ;
        RECT 4.000 356.640 495.600 358.040 ;
        RECT 4.000 354.640 496.000 356.640 ;
        RECT 4.400 353.240 495.600 354.640 ;
        RECT 4.000 351.240 496.000 353.240 ;
        RECT 4.400 349.840 495.600 351.240 ;
        RECT 4.000 347.840 496.000 349.840 ;
        RECT 4.400 346.440 495.600 347.840 ;
        RECT 4.000 344.440 496.000 346.440 ;
        RECT 4.400 343.040 495.600 344.440 ;
        RECT 4.000 341.040 496.000 343.040 ;
        RECT 4.400 339.640 495.600 341.040 ;
        RECT 4.000 337.640 496.000 339.640 ;
        RECT 4.400 336.240 495.600 337.640 ;
        RECT 4.000 334.240 496.000 336.240 ;
        RECT 4.400 332.840 496.000 334.240 ;
        RECT 4.000 330.840 496.000 332.840 ;
        RECT 4.400 329.440 495.600 330.840 ;
        RECT 4.000 327.440 496.000 329.440 ;
        RECT 4.400 326.040 495.600 327.440 ;
        RECT 4.000 324.040 496.000 326.040 ;
        RECT 4.400 322.640 495.600 324.040 ;
        RECT 4.000 320.640 496.000 322.640 ;
        RECT 4.400 319.240 495.600 320.640 ;
        RECT 4.000 317.240 496.000 319.240 ;
        RECT 4.400 315.840 495.600 317.240 ;
        RECT 4.000 313.840 496.000 315.840 ;
        RECT 4.000 312.440 495.600 313.840 ;
        RECT 4.000 310.440 496.000 312.440 ;
        RECT 4.400 309.040 495.600 310.440 ;
        RECT 4.000 307.040 496.000 309.040 ;
        RECT 4.400 305.640 495.600 307.040 ;
        RECT 4.000 303.640 496.000 305.640 ;
        RECT 4.400 302.240 495.600 303.640 ;
        RECT 4.000 300.240 496.000 302.240 ;
        RECT 4.400 298.840 495.600 300.240 ;
        RECT 4.000 296.840 496.000 298.840 ;
        RECT 4.400 295.440 495.600 296.840 ;
        RECT 4.000 293.440 496.000 295.440 ;
        RECT 4.400 292.040 495.600 293.440 ;
        RECT 4.000 290.040 496.000 292.040 ;
        RECT 4.400 288.640 495.600 290.040 ;
        RECT 4.000 286.640 496.000 288.640 ;
        RECT 4.400 285.240 496.000 286.640 ;
        RECT 4.000 283.240 496.000 285.240 ;
        RECT 4.400 281.840 495.600 283.240 ;
        RECT 4.000 279.840 496.000 281.840 ;
        RECT 4.400 278.440 495.600 279.840 ;
        RECT 4.000 276.440 496.000 278.440 ;
        RECT 4.400 275.040 495.600 276.440 ;
        RECT 4.000 273.040 496.000 275.040 ;
        RECT 4.400 271.640 495.600 273.040 ;
        RECT 4.000 269.640 496.000 271.640 ;
        RECT 4.000 268.240 495.600 269.640 ;
        RECT 4.000 266.240 496.000 268.240 ;
        RECT 4.400 264.840 495.600 266.240 ;
        RECT 4.000 262.840 496.000 264.840 ;
        RECT 4.400 261.440 495.600 262.840 ;
        RECT 4.000 259.440 496.000 261.440 ;
        RECT 4.400 258.040 495.600 259.440 ;
        RECT 4.000 256.040 496.000 258.040 ;
        RECT 4.400 254.640 495.600 256.040 ;
        RECT 4.000 252.640 496.000 254.640 ;
        RECT 4.400 251.240 495.600 252.640 ;
        RECT 4.000 249.240 496.000 251.240 ;
        RECT 4.400 247.840 495.600 249.240 ;
        RECT 4.000 245.840 496.000 247.840 ;
        RECT 4.400 244.440 495.600 245.840 ;
        RECT 4.000 242.440 496.000 244.440 ;
        RECT 4.400 241.040 496.000 242.440 ;
        RECT 4.000 239.040 496.000 241.040 ;
        RECT 4.400 237.640 495.600 239.040 ;
        RECT 4.000 235.640 496.000 237.640 ;
        RECT 4.400 234.240 495.600 235.640 ;
        RECT 4.000 232.240 496.000 234.240 ;
        RECT 4.400 230.840 495.600 232.240 ;
        RECT 4.000 228.840 496.000 230.840 ;
        RECT 4.400 227.440 495.600 228.840 ;
        RECT 4.000 225.440 496.000 227.440 ;
        RECT 4.000 224.040 495.600 225.440 ;
        RECT 4.000 222.040 496.000 224.040 ;
        RECT 4.400 220.640 495.600 222.040 ;
        RECT 4.000 218.640 496.000 220.640 ;
        RECT 4.400 217.240 495.600 218.640 ;
        RECT 4.000 215.240 496.000 217.240 ;
        RECT 4.400 213.840 495.600 215.240 ;
        RECT 4.000 211.840 496.000 213.840 ;
        RECT 4.400 210.440 495.600 211.840 ;
        RECT 4.000 208.440 496.000 210.440 ;
        RECT 4.400 207.040 495.600 208.440 ;
        RECT 4.000 205.040 496.000 207.040 ;
        RECT 4.400 203.640 495.600 205.040 ;
        RECT 4.000 201.640 496.000 203.640 ;
        RECT 4.400 200.240 495.600 201.640 ;
        RECT 4.000 198.240 496.000 200.240 ;
        RECT 4.400 196.840 496.000 198.240 ;
        RECT 4.000 194.840 496.000 196.840 ;
        RECT 4.400 193.440 495.600 194.840 ;
        RECT 4.000 191.440 496.000 193.440 ;
        RECT 4.400 190.040 495.600 191.440 ;
        RECT 4.000 188.040 496.000 190.040 ;
        RECT 4.400 186.640 495.600 188.040 ;
        RECT 4.000 184.640 496.000 186.640 ;
        RECT 4.400 183.240 495.600 184.640 ;
        RECT 4.000 181.240 496.000 183.240 ;
        RECT 4.000 179.840 495.600 181.240 ;
        RECT 4.000 177.840 496.000 179.840 ;
        RECT 4.400 176.440 495.600 177.840 ;
        RECT 4.000 174.440 496.000 176.440 ;
        RECT 4.400 173.040 495.600 174.440 ;
        RECT 4.000 171.040 496.000 173.040 ;
        RECT 4.400 169.640 495.600 171.040 ;
        RECT 4.000 167.640 496.000 169.640 ;
        RECT 4.400 166.240 495.600 167.640 ;
        RECT 4.000 164.240 496.000 166.240 ;
        RECT 4.400 162.840 495.600 164.240 ;
        RECT 4.000 160.840 496.000 162.840 ;
        RECT 4.400 159.440 495.600 160.840 ;
        RECT 4.000 157.440 496.000 159.440 ;
        RECT 4.400 156.040 495.600 157.440 ;
        RECT 4.000 154.040 496.000 156.040 ;
        RECT 4.400 152.640 496.000 154.040 ;
        RECT 4.000 150.640 496.000 152.640 ;
        RECT 4.400 149.240 495.600 150.640 ;
        RECT 4.000 147.240 496.000 149.240 ;
        RECT 4.400 145.840 495.600 147.240 ;
        RECT 4.000 143.840 496.000 145.840 ;
        RECT 4.400 142.440 495.600 143.840 ;
        RECT 4.000 140.440 496.000 142.440 ;
        RECT 4.400 139.040 495.600 140.440 ;
        RECT 4.000 137.040 496.000 139.040 ;
        RECT 4.000 135.640 495.600 137.040 ;
        RECT 4.000 133.640 496.000 135.640 ;
        RECT 4.400 132.240 495.600 133.640 ;
        RECT 4.000 130.240 496.000 132.240 ;
        RECT 4.400 128.840 495.600 130.240 ;
        RECT 4.000 126.840 496.000 128.840 ;
        RECT 4.400 125.440 495.600 126.840 ;
        RECT 4.000 123.440 496.000 125.440 ;
        RECT 4.400 122.040 495.600 123.440 ;
        RECT 4.000 120.040 496.000 122.040 ;
        RECT 4.400 118.640 495.600 120.040 ;
        RECT 4.000 116.640 496.000 118.640 ;
        RECT 4.400 115.240 495.600 116.640 ;
        RECT 4.000 113.240 496.000 115.240 ;
        RECT 4.400 111.840 495.600 113.240 ;
        RECT 4.000 109.840 496.000 111.840 ;
        RECT 4.400 108.440 496.000 109.840 ;
        RECT 4.000 106.440 496.000 108.440 ;
        RECT 4.400 105.040 495.600 106.440 ;
        RECT 4.000 103.040 496.000 105.040 ;
        RECT 4.400 101.640 495.600 103.040 ;
        RECT 4.000 99.640 496.000 101.640 ;
        RECT 4.400 98.240 495.600 99.640 ;
        RECT 4.000 96.240 496.000 98.240 ;
        RECT 4.400 94.840 495.600 96.240 ;
        RECT 4.000 92.840 496.000 94.840 ;
        RECT 4.000 91.440 495.600 92.840 ;
        RECT 4.000 89.440 496.000 91.440 ;
        RECT 4.400 88.040 495.600 89.440 ;
        RECT 4.000 86.040 496.000 88.040 ;
        RECT 4.400 84.640 495.600 86.040 ;
        RECT 4.000 82.640 496.000 84.640 ;
        RECT 4.400 81.240 495.600 82.640 ;
        RECT 4.000 79.240 496.000 81.240 ;
        RECT 4.400 77.840 495.600 79.240 ;
        RECT 4.000 75.840 496.000 77.840 ;
        RECT 4.400 74.440 495.600 75.840 ;
        RECT 4.000 72.440 496.000 74.440 ;
        RECT 4.400 71.040 495.600 72.440 ;
        RECT 4.000 69.040 496.000 71.040 ;
        RECT 4.400 67.640 495.600 69.040 ;
        RECT 4.000 65.640 496.000 67.640 ;
        RECT 4.400 64.240 496.000 65.640 ;
        RECT 4.000 62.240 496.000 64.240 ;
        RECT 4.400 60.840 495.600 62.240 ;
        RECT 4.000 58.840 496.000 60.840 ;
        RECT 4.400 57.440 495.600 58.840 ;
        RECT 4.000 55.440 496.000 57.440 ;
        RECT 4.400 54.040 495.600 55.440 ;
        RECT 4.000 52.040 496.000 54.040 ;
        RECT 4.400 50.640 495.600 52.040 ;
        RECT 4.000 48.640 496.000 50.640 ;
        RECT 4.000 47.240 495.600 48.640 ;
        RECT 4.000 45.240 496.000 47.240 ;
        RECT 4.400 43.840 495.600 45.240 ;
        RECT 4.000 41.840 496.000 43.840 ;
        RECT 4.400 40.440 495.600 41.840 ;
        RECT 4.000 38.440 496.000 40.440 ;
        RECT 4.400 37.040 495.600 38.440 ;
        RECT 4.000 35.040 496.000 37.040 ;
        RECT 4.400 33.640 495.600 35.040 ;
        RECT 4.000 31.640 496.000 33.640 ;
        RECT 4.400 30.240 495.600 31.640 ;
        RECT 4.000 28.240 496.000 30.240 ;
        RECT 4.400 26.840 495.600 28.240 ;
        RECT 4.000 24.840 496.000 26.840 ;
        RECT 4.400 23.440 495.600 24.840 ;
        RECT 4.000 21.440 496.000 23.440 ;
        RECT 4.400 20.040 496.000 21.440 ;
        RECT 4.000 18.040 496.000 20.040 ;
        RECT 4.400 16.640 495.600 18.040 ;
        RECT 4.000 14.640 496.000 16.640 ;
        RECT 4.400 13.240 495.600 14.640 ;
        RECT 4.000 11.240 496.000 13.240 ;
        RECT 4.400 9.840 495.600 11.240 ;
        RECT 4.000 7.840 496.000 9.840 ;
        RECT 4.400 6.440 495.600 7.840 ;
        RECT 4.000 4.440 496.000 6.440 ;
        RECT 4.000 3.575 495.600 4.440 ;
      LAYER met4 ;
        RECT 244.095 12.415 244.425 414.625 ;
  END
END openram_testchip
END LIBRARY

