magic
tech sky130A
timestamp 1640667123
<< metal3 >>
rect -8417 249 -5118 1077
<< mimcap >>
rect -8361 1035 -5161 1063
rect -8361 1000 -8333 1035
rect -8298 1034 -5161 1035
rect -8298 1031 -7303 1034
rect -8298 1000 -7888 1031
rect -8361 996 -7888 1000
rect -7853 999 -7303 1031
rect -7268 1033 -5161 1034
rect -7268 999 -6708 1033
rect -7853 998 -6708 999
rect -6673 998 -6042 1033
rect -6007 998 -5273 1033
rect -5238 998 -5161 1033
rect -7853 996 -5161 998
rect -8361 321 -5161 996
rect -8361 318 -6105 321
rect -8361 283 -8341 318
rect -8306 283 -7852 318
rect -7817 283 -7287 318
rect -7252 317 -6105 318
rect -7252 283 -6748 317
rect -8361 282 -6748 283
rect -6713 286 -6105 317
rect -6070 317 -5161 321
rect -6070 286 -5279 317
rect -6713 282 -5279 286
rect -5244 282 -5161 317
rect -8361 263 -5161 282
<< mimcapcontact >>
rect -8333 1000 -8298 1035
rect -7888 996 -7853 1031
rect -7303 999 -7268 1034
rect -6708 998 -6673 1033
rect -6042 998 -6007 1033
rect -5273 998 -5238 1033
rect -8341 283 -8306 318
rect -7852 283 -7817 318
rect -7287 283 -7252 318
rect -6748 282 -6713 317
rect -6105 286 -6070 321
rect -5279 282 -5244 317
<< metal4 >>
rect -8345 1035 -5177 1045
rect -8345 1000 -8333 1035
rect -8298 1034 -5177 1035
rect -8298 1031 -7303 1034
rect -8298 1000 -7888 1031
rect -8345 996 -7888 1000
rect -7853 999 -7303 1031
rect -7268 1033 -5177 1034
rect -7268 999 -6708 1033
rect -7853 998 -6708 999
rect -6673 998 -6042 1033
rect -6007 998 -5273 1033
rect -5238 998 -5177 1033
rect -7853 996 -5177 998
rect -8345 990 -5177 996
rect -8349 321 -5181 328
rect -8349 318 -6105 321
rect -8349 283 -8341 318
rect -8306 283 -7852 318
rect -7817 283 -7287 318
rect -7252 317 -6105 318
rect -7252 283 -6748 317
rect -8349 282 -6748 283
rect -6713 286 -6105 317
rect -6070 317 -5181 321
rect -6070 286 -5279 317
rect -6713 282 -5279 286
rect -5244 282 -5181 317
rect -8349 273 -5181 282
<< end >>
