VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_32_512_sky130
   CLASS BLOCK ;
   SIZE 475.02 BY 319.3 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.56 0.0 113.94 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.0 0.0 119.38 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.12 0.0 125.5 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 0.0 130.94 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.68 0.0 137.06 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.48 0.0 143.86 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.36 0.0 154.74 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 0.0 160.18 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 0.0 166.3 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.36 0.0 171.74 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.48 0.0 177.86 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.6 0.0 183.98 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 0.0 189.42 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.84 0.0 196.22 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 0.0 207.78 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.52 0.0 213.9 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.28 0.0 218.66 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  225.08 0.0 225.46 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  236.64 0.0 237.02 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 0.0 243.14 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 0.0 248.58 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 0.0 260.14 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 0.0 271.7 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.76 0.0 277.14 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.88 0.0 283.26 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  295.12 0.0 295.5 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  299.88 0.0 300.26 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.2 0.0 78.58 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.32 0.0 84.7 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.72 0.38 139.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 147.56 0.38 147.94 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 152.32 0.38 152.7 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.2 0.38 163.58 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.96 0.38 168.34 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 175.44 0.38 175.82 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 181.56 0.38 181.94 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.72 0.38 37.1 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 43.52 0.38 43.9 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 37.4 0.38 37.78 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  90.44 0.0 90.82 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.88 0.0 96.26 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.68 0.0 103.06 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.12 0.0 108.5 0.38 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  306.68 0.0 307.06 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 0.0 140.46 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 0.0 152.02 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.04 0.0 172.42 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  181.56 0.0 181.94 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 0.0 192.14 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  201.96 0.0 202.34 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.8 0.0 211.18 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.32 0.0 220.7 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 0.0 232.26 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.08 0.0 242.46 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  251.6 0.0 251.98 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  261.8 0.0 262.18 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 0.0 272.38 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 0.0 281.22 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.72 0.0 292.1 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 0.0 300.94 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 0.0 310.46 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 0.0 322.02 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.84 0.0 332.22 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  351.56 0.0 351.94 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.76 0.0 362.14 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 0.0 372.34 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  380.12 0.0 380.5 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  391.68 0.0 392.06 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  401.88 0.0 402.26 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  411.4 0.0 411.78 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  474.64 58.48 475.02 58.86 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  474.64 59.16 475.02 59.54 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  474.64 63.92 475.02 64.3 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  474.64 59.84 475.02 60.22 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  474.64 61.88 475.02 62.26 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  1.36 317.56 473.66 319.3 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 319.3 ;
         LAYER met3 ;
         RECT  1.36 1.36 473.66 3.1 ;
         LAYER met4 ;
         RECT  471.92 1.36 473.66 319.3 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 470.26 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 315.9 ;
         LAYER met3 ;
         RECT  4.76 314.16 470.26 315.9 ;
         LAYER met4 ;
         RECT  468.52 4.76 470.26 315.9 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 474.4 318.68 ;
   LAYER  met2 ;
      RECT  0.62 0.62 474.4 318.68 ;
   LAYER  met3 ;
      RECT  0.98 138.12 474.4 139.7 ;
      RECT  0.62 139.7 0.98 146.96 ;
      RECT  0.62 148.54 0.98 151.72 ;
      RECT  0.62 153.3 0.98 162.6 ;
      RECT  0.62 164.18 0.98 167.36 ;
      RECT  0.62 168.94 0.98 174.84 ;
      RECT  0.62 176.42 0.98 180.96 ;
      RECT  0.62 44.5 0.98 138.12 ;
      RECT  0.62 38.38 0.98 42.92 ;
      RECT  0.98 57.88 474.04 59.46 ;
      RECT  0.98 59.46 474.04 138.12 ;
      RECT  474.04 64.9 474.4 138.12 ;
      RECT  474.04 60.82 474.4 61.28 ;
      RECT  474.04 62.86 474.4 63.32 ;
      RECT  474.26 139.7 474.4 316.96 ;
      RECT  474.26 316.96 474.4 318.68 ;
      RECT  0.62 182.54 0.76 316.96 ;
      RECT  0.62 316.96 0.76 318.68 ;
      RECT  0.76 182.54 0.98 316.96 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 36.12 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 36.12 ;
      RECT  0.98 0.62 474.04 0.76 ;
      RECT  474.04 0.62 474.26 0.76 ;
      RECT  474.04 3.7 474.26 57.88 ;
      RECT  474.26 0.62 474.4 0.76 ;
      RECT  474.26 0.76 474.4 3.7 ;
      RECT  474.26 3.7 474.4 57.88 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 57.88 ;
      RECT  4.16 3.7 470.86 4.16 ;
      RECT  4.16 7.1 470.86 57.88 ;
      RECT  470.86 3.7 474.04 4.16 ;
      RECT  470.86 4.16 474.04 7.1 ;
      RECT  470.86 7.1 474.04 57.88 ;
      RECT  0.98 139.7 4.16 313.56 ;
      RECT  0.98 313.56 4.16 316.5 ;
      RECT  0.98 316.5 4.16 316.96 ;
      RECT  4.16 139.7 470.86 313.56 ;
      RECT  4.16 316.5 470.86 316.96 ;
      RECT  470.86 139.7 474.26 313.56 ;
      RECT  470.86 313.56 474.26 316.5 ;
      RECT  470.86 316.5 474.26 316.96 ;
   LAYER  met4 ;
      RECT  112.96 0.98 114.54 318.68 ;
      RECT  114.54 0.62 118.4 0.98 ;
      RECT  119.98 0.62 124.52 0.98 ;
      RECT  126.1 0.62 129.96 0.98 ;
      RECT  131.54 0.62 136.08 0.98 ;
      RECT  144.46 0.62 147.64 0.98 ;
      RECT  155.34 0.62 159.2 0.98 ;
      RECT  166.9 0.62 170.76 0.98 ;
      RECT  184.58 0.62 188.44 0.98 ;
      RECT  196.82 0.62 200.68 0.98 ;
      RECT  214.5 0.62 217.68 0.98 ;
      RECT  226.06 0.62 229.92 0.98 ;
      RECT  243.74 0.62 247.6 0.98 ;
      RECT  254.62 0.62 259.16 0.98 ;
      RECT  266.86 0.62 270.72 0.98 ;
      RECT  283.86 0.62 287.72 0.98 ;
      RECT  296.1 0.62 299.28 0.98 ;
      RECT  79.18 0.62 83.72 0.98 ;
      RECT  85.3 0.62 89.84 0.98 ;
      RECT  91.42 0.62 95.28 0.98 ;
      RECT  96.86 0.62 102.08 0.98 ;
      RECT  103.66 0.62 107.52 0.98 ;
      RECT  109.1 0.62 112.96 0.98 ;
      RECT  137.66 0.62 139.48 0.98 ;
      RECT  141.06 0.62 142.88 0.98 ;
      RECT  149.22 0.62 151.04 0.98 ;
      RECT  152.62 0.62 153.76 0.98 ;
      RECT  160.78 0.62 161.24 0.98 ;
      RECT  162.82 0.62 165.32 0.98 ;
      RECT  173.02 0.62 176.88 0.98 ;
      RECT  178.46 0.62 180.96 0.98 ;
      RECT  182.54 0.62 183.0 0.98 ;
      RECT  190.02 0.62 191.16 0.98 ;
      RECT  192.74 0.62 195.24 0.98 ;
      RECT  202.94 0.62 206.8 0.98 ;
      RECT  208.38 0.62 210.2 0.98 ;
      RECT  211.78 0.62 212.92 0.98 ;
      RECT  219.26 0.62 219.72 0.98 ;
      RECT  221.3 0.62 224.48 0.98 ;
      RECT  232.86 0.62 236.04 0.98 ;
      RECT  237.62 0.62 241.48 0.98 ;
      RECT  249.18 0.62 251.0 0.98 ;
      RECT  252.58 0.62 253.04 0.98 ;
      RECT  260.74 0.62 261.2 0.98 ;
      RECT  262.78 0.62 265.28 0.98 ;
      RECT  272.98 0.62 276.16 0.98 ;
      RECT  277.74 0.62 280.24 0.98 ;
      RECT  281.82 0.62 282.28 0.98 ;
      RECT  289.3 0.62 291.12 0.98 ;
      RECT  292.7 0.62 294.52 0.98 ;
      RECT  301.54 0.62 306.08 0.98 ;
      RECT  307.66 0.62 309.48 0.98 ;
      RECT  311.06 0.62 321.04 0.98 ;
      RECT  322.62 0.62 331.24 0.98 ;
      RECT  332.82 0.62 340.76 0.98 ;
      RECT  342.34 0.62 350.96 0.98 ;
      RECT  352.54 0.62 361.16 0.98 ;
      RECT  362.74 0.62 371.36 0.98 ;
      RECT  372.94 0.62 379.52 0.98 ;
      RECT  381.1 0.62 391.08 0.98 ;
      RECT  392.66 0.62 401.28 0.98 ;
      RECT  402.86 0.62 410.8 0.98 ;
      RECT  0.62 0.98 0.76 318.68 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 77.6 0.76 ;
      RECT  3.7 0.76 77.6 0.98 ;
      RECT  474.26 0.98 474.4 318.68 ;
      RECT  412.38 0.62 471.32 0.76 ;
      RECT  412.38 0.76 471.32 0.98 ;
      RECT  471.32 0.62 474.26 0.76 ;
      RECT  474.26 0.62 474.4 0.76 ;
      RECT  474.26 0.76 474.4 0.98 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 316.5 ;
      RECT  3.7 316.5 4.16 318.68 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 316.5 7.1 318.68 ;
      RECT  7.1 0.98 112.96 4.16 ;
      RECT  7.1 4.16 112.96 316.5 ;
      RECT  7.1 316.5 112.96 318.68 ;
      RECT  114.54 0.98 467.92 4.16 ;
      RECT  114.54 4.16 467.92 316.5 ;
      RECT  114.54 316.5 467.92 318.68 ;
      RECT  467.92 0.98 470.86 4.16 ;
      RECT  467.92 316.5 470.86 318.68 ;
      RECT  470.86 0.98 471.32 4.16 ;
      RECT  470.86 4.16 471.32 316.5 ;
      RECT  470.86 316.5 471.32 318.68 ;
   END
END    sram_1rw0r0w_32_512_sky130
END    LIBRARY
