// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

`timescale 1 ns / 1 ps

module io_ports_tb;
	reg clock;
	reg RSTB;
	reg CSB;
	reg power1, power2;
	reg power3, power4;

	wire gpio;
	wire [37:0] mprj_io;
	wire [37:0] mprj_io_0;

	assign mprj_io_0 = mprj_io[37:0];
	// assign mprj_io_0 = {mprj_io[8:4],mprj_io[2:0]};

	assign mprj_io[3] = (CSB == 1'b1) ? 1'b1 : 1'bz;
	// assign mprj_io[3] = 1'b1;

	// External clock is used by default.  Make this artificially fast for the
	// simulation.  Normally this would be a slow clock and the digital PLL
	// would be the fast clock.

	always #12.5 clock <= (clock === 1'b0);

	initial begin
		clock = 0;
	end

	initial begin
		$dumpfile("io_ports.vcd");
		$dumpvars(0, io_ports_tb);

		// Repeat cycles of 10000 clock edges as needed to complete testbench
		repeat (25) begin
			repeat (10000	) @(posedge clock);
			// $display("+10000 cycles");
		end
		$display("%c[1;31m",27);
		`ifdef GL
			$display ("Monitor: Timeout, Test Mega-Project IO Ports (GL) Failed");
		`else
			$display ("Monitor: Timeout, Test Mega-Project IO Ports (RTL) Failed");
		`endif
		$display("%c[0m",27);
		$finish;
	end

	initial begin
	    // Observe Output pins
		wait(mprj_io_0 == 38'h0000000001);
		wait(mprj_io_0 == 38'h2000000000);
		wait(mprj_io_0 == 38'h3000000000);
		wait(mprj_io_0 == 38'h3800000000);
		wait(mprj_io_0 == 38'h3C00000000);
		wait(mprj_io_0 == 38'h3E00000000);
		wait(mprj_io_0 == 38'h3F00000000);
		wait(mprj_io_0 == 38'h3F80000000);
		wait(mprj_io_0 == 38'h3FC0000000);
		wait(mprj_io_0 == 38'h3FE0000000);
		wait(mprj_io_0 == 38'h3FF0000000);
		wait(mprj_io_0 == 38'h3FF8000000);
		wait(mprj_io_0 == 38'h3FFC000000);
		wait(mprj_io_0 == 38'h3FFE000000);
		wait(mprj_io_0 == 38'h3FFF000000);
		wait(mprj_io_0 == 38'h3FFF800000);
		wait(mprj_io_0 == 38'h3FFFC00000);
		wait(mprj_io_0 == 38'h3FFFE00000);
		wait(mprj_io_0 == 38'h3FFFF00000);
		wait(mprj_io_0 == 38'h3FFFF80000);
		wait(mprj_io_0 == 38'h3FFFFC0000);
		wait(mprj_io_0 == 38'h3FFFFE0000);
		wait(mprj_io_0 == 38'h3FFFFF0000);
		wait(mprj_io_0 == 38'h3FFFFF8000);
		wait(mprj_io_0 == 38'h3FFFFFC000);
		wait(mprj_io_0 == 38'h3FFFFFE000);
		wait(mprj_io_0 == 38'h3FFFFFF000);
		wait(mprj_io_0 == 38'h3FFFFFF800);
		wait(mprj_io_0 == 38'h3FFFFFFC00);
		wait(mprj_io_0 == 38'h3FFFFFFE00);
		wait(mprj_io_0 == 38'h3FFFFFFF00);
		wait(mprj_io_0 == 38'h3FFFFFFF80);
		wait(mprj_io_0 == 38'h3FFFFFFFC0);
		wait(mprj_io_0 == 38'h3FFFFFFFE0);
		wait(mprj_io_0 == 38'h3FFFFFFFF0);
		wait(mprj_io_0 == 38'h3FFFFFFFF8);
		wait(mprj_io_0 == 38'h3FFFFFFFFC);
		wait(mprj_io_0 == 38'h3FFFFFFFFE);
		wait(mprj_io_0 == 38'h3FFFFFFFFF);
		wait(mprj_io_0 == 38'h0000000000);
		
		`ifdef GL
	    	$display("Monitor: Test 1 Mega-Project IO (GL) Passed");
		`else
		    $display("Monitor: Test 1 Mega-Project IO (RTL) Passed");
		`endif
	    $finish;
	end

	initial begin
		RSTB <= 1'b0;
		CSB  <= 1'b1;		// Force CSB high
		#2000;
		RSTB <= 1'b1;	    	// Release reset
		#300000;
		CSB = 1'b0;		// CSB can be released
	end

	initial begin		// Power-up sequence
		power1 <= 1'b0;
		power2 <= 1'b0;
		power3 <= 1'b0;
		power4 <= 1'b0;
		#100;
		power1 <= 1'b1;
		#100;
		power2 <= 1'b1;
		#100;
		power3 <= 1'b1;
		#100;
		power4 <= 1'b1;
	end

	always @(mprj_io) begin
		#1 $display("MPRJ-IO state = %b ", mprj_io[37:0]);
	end

	wire flash_csb;
	wire flash_clk;
	wire flash_io0;
	wire flash_io1;

	wire VDD3V3;
	wire VDD1V8;
	wire VSS;
	
	assign VDD3V3 = power1;
	assign VDD1V8 = power2;
	assign VSS = 1'b0;

	caravel uut (
		.vddio	  (VDD3V3),
		.vddio_2  (VDD3V3),
		.vssio	  (VSS),
		.vssio_2  (VSS),
		.vdda	  (VDD3V3),
		.vssa	  (VSS),
		.vccd	  (VDD1V8),
		.vssd	  (VSS),
		.vdda1    (VDD3V3),
		.vdda1_2  (VDD3V3),
		.vdda2    (VDD3V3),
		.vssa1	  (VSS),
		.vssa1_2  (VSS),
		.vssa2	  (VSS),
		.vccd1	  (VDD1V8),
		.vccd2	  (VDD1V8),
		.vssd1	  (VSS),
		.vssd2	  (VSS),
		.clock    (clock),
		.gpio     (gpio),
		.mprj_io  (mprj_io),
		.flash_csb(flash_csb),
		.flash_clk(flash_clk),
		.flash_io0(flash_io0),
		.flash_io1(flash_io1),
		.resetb	  (RSTB)
	);

	spiflash #(
		.FILENAME("io_ports.hex")
	) spiflash (
		.csb(flash_csb),
		.clk(flash_clk),
		.io0(flash_io0),
		.io1(flash_io1),
		.io2(),			// not used
		.io3()			// not used
	);

endmodule
`default_nettype wire
