magic
tech sky130A
magscale 1 2
timestamp 1624051196
<< obsli1 >>
rect 1104 1853 582820 701777
<< obsm1 >>
rect 1104 1572 583450 701808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 1674 703464 8030 703520
rect 8254 703464 24222 703520
rect 24446 703464 40414 703520
rect 40638 703464 56698 703520
rect 56922 703464 72890 703520
rect 73114 703464 89082 703520
rect 89306 703464 105366 703520
rect 105590 703464 121558 703520
rect 121782 703464 137750 703520
rect 137974 703464 154034 703520
rect 154258 703464 170226 703520
rect 170450 703464 186418 703520
rect 186642 703464 202702 703520
rect 202926 703464 218894 703520
rect 219118 703464 235086 703520
rect 235310 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 300038 703520
rect 300262 703464 316230 703520
rect 316454 703464 332422 703520
rect 332646 703464 348706 703520
rect 348930 703464 364898 703520
rect 365122 703464 381090 703520
rect 381314 703464 397374 703520
rect 397598 703464 413566 703520
rect 413790 703464 429758 703520
rect 429982 703464 446042 703520
rect 446266 703464 462234 703520
rect 462458 703464 478426 703520
rect 478650 703464 494710 703520
rect 494934 703464 510902 703520
rect 511126 703464 527094 703520
rect 527318 703464 543378 703520
rect 543602 703464 559570 703520
rect 559794 703464 575762 703520
rect 575986 703464 583444 703520
rect 1674 536 583444 703464
rect 1814 480 2786 536
rect 3010 480 3982 536
rect 4206 480 5178 536
rect 5402 480 6374 536
rect 6598 480 7570 536
rect 7794 480 8674 536
rect 8898 480 9870 536
rect 10094 480 11066 536
rect 11290 480 12262 536
rect 12486 480 13458 536
rect 13682 480 14654 536
rect 14878 480 15850 536
rect 16074 480 16954 536
rect 17178 480 18150 536
rect 18374 480 19346 536
rect 19570 480 20542 536
rect 20766 480 21738 536
rect 21962 480 22934 536
rect 23158 480 24130 536
rect 24354 480 25234 536
rect 25458 480 26430 536
rect 26654 480 27626 536
rect 27850 480 28822 536
rect 29046 480 30018 536
rect 30242 480 31214 536
rect 31438 480 32318 536
rect 32542 480 33514 536
rect 33738 480 34710 536
rect 34934 480 35906 536
rect 36130 480 37102 536
rect 37326 480 38298 536
rect 38522 480 39494 536
rect 39718 480 40598 536
rect 40822 480 41794 536
rect 42018 480 42990 536
rect 43214 480 44186 536
rect 44410 480 45382 536
rect 45606 480 46578 536
rect 46802 480 47774 536
rect 47998 480 48878 536
rect 49102 480 50074 536
rect 50298 480 51270 536
rect 51494 480 52466 536
rect 52690 480 53662 536
rect 53886 480 54858 536
rect 55082 480 55962 536
rect 56186 480 57158 536
rect 57382 480 58354 536
rect 58578 480 59550 536
rect 59774 480 60746 536
rect 60970 480 61942 536
rect 62166 480 63138 536
rect 63362 480 64242 536
rect 64466 480 65438 536
rect 65662 480 66634 536
rect 66858 480 67830 536
rect 68054 480 69026 536
rect 69250 480 70222 536
rect 70446 480 71418 536
rect 71642 480 72522 536
rect 72746 480 73718 536
rect 73942 480 74914 536
rect 75138 480 76110 536
rect 76334 480 77306 536
rect 77530 480 78502 536
rect 78726 480 79606 536
rect 79830 480 80802 536
rect 81026 480 81998 536
rect 82222 480 83194 536
rect 83418 480 84390 536
rect 84614 480 85586 536
rect 85810 480 86782 536
rect 87006 480 87886 536
rect 88110 480 89082 536
rect 89306 480 90278 536
rect 90502 480 91474 536
rect 91698 480 92670 536
rect 92894 480 93866 536
rect 94090 480 95062 536
rect 95286 480 96166 536
rect 96390 480 97362 536
rect 97586 480 98558 536
rect 98782 480 99754 536
rect 99978 480 100950 536
rect 101174 480 102146 536
rect 102370 480 103250 536
rect 103474 480 104446 536
rect 104670 480 105642 536
rect 105866 480 106838 536
rect 107062 480 108034 536
rect 108258 480 109230 536
rect 109454 480 110426 536
rect 110650 480 111530 536
rect 111754 480 112726 536
rect 112950 480 113922 536
rect 114146 480 115118 536
rect 115342 480 116314 536
rect 116538 480 117510 536
rect 117734 480 118706 536
rect 118930 480 119810 536
rect 120034 480 121006 536
rect 121230 480 122202 536
rect 122426 480 123398 536
rect 123622 480 124594 536
rect 124818 480 125790 536
rect 126014 480 126894 536
rect 127118 480 128090 536
rect 128314 480 129286 536
rect 129510 480 130482 536
rect 130706 480 131678 536
rect 131902 480 132874 536
rect 133098 480 134070 536
rect 134294 480 135174 536
rect 135398 480 136370 536
rect 136594 480 137566 536
rect 137790 480 138762 536
rect 138986 480 139958 536
rect 140182 480 141154 536
rect 141378 480 142350 536
rect 142574 480 143454 536
rect 143678 480 144650 536
rect 144874 480 145846 536
rect 146070 480 147042 536
rect 147266 480 148238 536
rect 148462 480 149434 536
rect 149658 480 150538 536
rect 150762 480 151734 536
rect 151958 480 152930 536
rect 153154 480 154126 536
rect 154350 480 155322 536
rect 155546 480 156518 536
rect 156742 480 157714 536
rect 157938 480 158818 536
rect 159042 480 160014 536
rect 160238 480 161210 536
rect 161434 480 162406 536
rect 162630 480 163602 536
rect 163826 480 164798 536
rect 165022 480 165994 536
rect 166218 480 167098 536
rect 167322 480 168294 536
rect 168518 480 169490 536
rect 169714 480 170686 536
rect 170910 480 171882 536
rect 172106 480 173078 536
rect 173302 480 174182 536
rect 174406 480 175378 536
rect 175602 480 176574 536
rect 176798 480 177770 536
rect 177994 480 178966 536
rect 179190 480 180162 536
rect 180386 480 181358 536
rect 181582 480 182462 536
rect 182686 480 183658 536
rect 183882 480 184854 536
rect 185078 480 186050 536
rect 186274 480 187246 536
rect 187470 480 188442 536
rect 188666 480 189638 536
rect 189862 480 190742 536
rect 190966 480 191938 536
rect 192162 480 193134 536
rect 193358 480 194330 536
rect 194554 480 195526 536
rect 195750 480 196722 536
rect 196946 480 197826 536
rect 198050 480 199022 536
rect 199246 480 200218 536
rect 200442 480 201414 536
rect 201638 480 202610 536
rect 202834 480 203806 536
rect 204030 480 205002 536
rect 205226 480 206106 536
rect 206330 480 207302 536
rect 207526 480 208498 536
rect 208722 480 209694 536
rect 209918 480 210890 536
rect 211114 480 212086 536
rect 212310 480 213282 536
rect 213506 480 214386 536
rect 214610 480 215582 536
rect 215806 480 216778 536
rect 217002 480 217974 536
rect 218198 480 219170 536
rect 219394 480 220366 536
rect 220590 480 221470 536
rect 221694 480 222666 536
rect 222890 480 223862 536
rect 224086 480 225058 536
rect 225282 480 226254 536
rect 226478 480 227450 536
rect 227674 480 228646 536
rect 228870 480 229750 536
rect 229974 480 230946 536
rect 231170 480 232142 536
rect 232366 480 233338 536
rect 233562 480 234534 536
rect 234758 480 235730 536
rect 235954 480 236926 536
rect 237150 480 238030 536
rect 238254 480 239226 536
rect 239450 480 240422 536
rect 240646 480 241618 536
rect 241842 480 242814 536
rect 243038 480 244010 536
rect 244234 480 245114 536
rect 245338 480 246310 536
rect 246534 480 247506 536
rect 247730 480 248702 536
rect 248926 480 249898 536
rect 250122 480 251094 536
rect 251318 480 252290 536
rect 252514 480 253394 536
rect 253618 480 254590 536
rect 254814 480 255786 536
rect 256010 480 256982 536
rect 257206 480 258178 536
rect 258402 480 259374 536
rect 259598 480 260570 536
rect 260794 480 261674 536
rect 261898 480 262870 536
rect 263094 480 264066 536
rect 264290 480 265262 536
rect 265486 480 266458 536
rect 266682 480 267654 536
rect 267878 480 268758 536
rect 268982 480 269954 536
rect 270178 480 271150 536
rect 271374 480 272346 536
rect 272570 480 273542 536
rect 273766 480 274738 536
rect 274962 480 275934 536
rect 276158 480 277038 536
rect 277262 480 278234 536
rect 278458 480 279430 536
rect 279654 480 280626 536
rect 280850 480 281822 536
rect 282046 480 283018 536
rect 283242 480 284214 536
rect 284438 480 285318 536
rect 285542 480 286514 536
rect 286738 480 287710 536
rect 287934 480 288906 536
rect 289130 480 290102 536
rect 290326 480 291298 536
rect 291522 480 292494 536
rect 292718 480 293598 536
rect 293822 480 294794 536
rect 295018 480 295990 536
rect 296214 480 297186 536
rect 297410 480 298382 536
rect 298606 480 299578 536
rect 299802 480 300682 536
rect 300906 480 301878 536
rect 302102 480 303074 536
rect 303298 480 304270 536
rect 304494 480 305466 536
rect 305690 480 306662 536
rect 306886 480 307858 536
rect 308082 480 308962 536
rect 309186 480 310158 536
rect 310382 480 311354 536
rect 311578 480 312550 536
rect 312774 480 313746 536
rect 313970 480 314942 536
rect 315166 480 316138 536
rect 316362 480 317242 536
rect 317466 480 318438 536
rect 318662 480 319634 536
rect 319858 480 320830 536
rect 321054 480 322026 536
rect 322250 480 323222 536
rect 323446 480 324326 536
rect 324550 480 325522 536
rect 325746 480 326718 536
rect 326942 480 327914 536
rect 328138 480 329110 536
rect 329334 480 330306 536
rect 330530 480 331502 536
rect 331726 480 332606 536
rect 332830 480 333802 536
rect 334026 480 334998 536
rect 335222 480 336194 536
rect 336418 480 337390 536
rect 337614 480 338586 536
rect 338810 480 339782 536
rect 340006 480 340886 536
rect 341110 480 342082 536
rect 342306 480 343278 536
rect 343502 480 344474 536
rect 344698 480 345670 536
rect 345894 480 346866 536
rect 347090 480 347970 536
rect 348194 480 349166 536
rect 349390 480 350362 536
rect 350586 480 351558 536
rect 351782 480 352754 536
rect 352978 480 353950 536
rect 354174 480 355146 536
rect 355370 480 356250 536
rect 356474 480 357446 536
rect 357670 480 358642 536
rect 358866 480 359838 536
rect 360062 480 361034 536
rect 361258 480 362230 536
rect 362454 480 363426 536
rect 363650 480 364530 536
rect 364754 480 365726 536
rect 365950 480 366922 536
rect 367146 480 368118 536
rect 368342 480 369314 536
rect 369538 480 370510 536
rect 370734 480 371614 536
rect 371838 480 372810 536
rect 373034 480 374006 536
rect 374230 480 375202 536
rect 375426 480 376398 536
rect 376622 480 377594 536
rect 377818 480 378790 536
rect 379014 480 379894 536
rect 380118 480 381090 536
rect 381314 480 382286 536
rect 382510 480 383482 536
rect 383706 480 384678 536
rect 384902 480 385874 536
rect 386098 480 387070 536
rect 387294 480 388174 536
rect 388398 480 389370 536
rect 389594 480 390566 536
rect 390790 480 391762 536
rect 391986 480 392958 536
rect 393182 480 394154 536
rect 394378 480 395258 536
rect 395482 480 396454 536
rect 396678 480 397650 536
rect 397874 480 398846 536
rect 399070 480 400042 536
rect 400266 480 401238 536
rect 401462 480 402434 536
rect 402658 480 403538 536
rect 403762 480 404734 536
rect 404958 480 405930 536
rect 406154 480 407126 536
rect 407350 480 408322 536
rect 408546 480 409518 536
rect 409742 480 410714 536
rect 410938 480 411818 536
rect 412042 480 413014 536
rect 413238 480 414210 536
rect 414434 480 415406 536
rect 415630 480 416602 536
rect 416826 480 417798 536
rect 418022 480 418902 536
rect 419126 480 420098 536
rect 420322 480 421294 536
rect 421518 480 422490 536
rect 422714 480 423686 536
rect 423910 480 424882 536
rect 425106 480 426078 536
rect 426302 480 427182 536
rect 427406 480 428378 536
rect 428602 480 429574 536
rect 429798 480 430770 536
rect 430994 480 431966 536
rect 432190 480 433162 536
rect 433386 480 434358 536
rect 434582 480 435462 536
rect 435686 480 436658 536
rect 436882 480 437854 536
rect 438078 480 439050 536
rect 439274 480 440246 536
rect 440470 480 441442 536
rect 441666 480 442546 536
rect 442770 480 443742 536
rect 443966 480 444938 536
rect 445162 480 446134 536
rect 446358 480 447330 536
rect 447554 480 448526 536
rect 448750 480 449722 536
rect 449946 480 450826 536
rect 451050 480 452022 536
rect 452246 480 453218 536
rect 453442 480 454414 536
rect 454638 480 455610 536
rect 455834 480 456806 536
rect 457030 480 458002 536
rect 458226 480 459106 536
rect 459330 480 460302 536
rect 460526 480 461498 536
rect 461722 480 462694 536
rect 462918 480 463890 536
rect 464114 480 465086 536
rect 465310 480 466190 536
rect 466414 480 467386 536
rect 467610 480 468582 536
rect 468806 480 469778 536
rect 470002 480 470974 536
rect 471198 480 472170 536
rect 472394 480 473366 536
rect 473590 480 474470 536
rect 474694 480 475666 536
rect 475890 480 476862 536
rect 477086 480 478058 536
rect 478282 480 479254 536
rect 479478 480 480450 536
rect 480674 480 481646 536
rect 481870 480 482750 536
rect 482974 480 483946 536
rect 484170 480 485142 536
rect 485366 480 486338 536
rect 486562 480 487534 536
rect 487758 480 488730 536
rect 488954 480 489834 536
rect 490058 480 491030 536
rect 491254 480 492226 536
rect 492450 480 493422 536
rect 493646 480 494618 536
rect 494842 480 495814 536
rect 496038 480 497010 536
rect 497234 480 498114 536
rect 498338 480 499310 536
rect 499534 480 500506 536
rect 500730 480 501702 536
rect 501926 480 502898 536
rect 503122 480 504094 536
rect 504318 480 505290 536
rect 505514 480 506394 536
rect 506618 480 507590 536
rect 507814 480 508786 536
rect 509010 480 509982 536
rect 510206 480 511178 536
rect 511402 480 512374 536
rect 512598 480 513478 536
rect 513702 480 514674 536
rect 514898 480 515870 536
rect 516094 480 517066 536
rect 517290 480 518262 536
rect 518486 480 519458 536
rect 519682 480 520654 536
rect 520878 480 521758 536
rect 521982 480 522954 536
rect 523178 480 524150 536
rect 524374 480 525346 536
rect 525570 480 526542 536
rect 526766 480 527738 536
rect 527962 480 528934 536
rect 529158 480 530038 536
rect 530262 480 531234 536
rect 531458 480 532430 536
rect 532654 480 533626 536
rect 533850 480 534822 536
rect 535046 480 536018 536
rect 536242 480 537122 536
rect 537346 480 538318 536
rect 538542 480 539514 536
rect 539738 480 540710 536
rect 540934 480 541906 536
rect 542130 480 543102 536
rect 543326 480 544298 536
rect 544522 480 545402 536
rect 545626 480 546598 536
rect 546822 480 547794 536
rect 548018 480 548990 536
rect 549214 480 550186 536
rect 550410 480 551382 536
rect 551606 480 552578 536
rect 552802 480 553682 536
rect 553906 480 554878 536
rect 555102 480 556074 536
rect 556298 480 557270 536
rect 557494 480 558466 536
rect 558690 480 559662 536
rect 559886 480 560766 536
rect 560990 480 561962 536
rect 562186 480 563158 536
rect 563382 480 564354 536
rect 564578 480 565550 536
rect 565774 480 566746 536
rect 566970 480 567942 536
rect 568166 480 569046 536
rect 569270 480 570242 536
rect 570466 480 571438 536
rect 571662 480 572634 536
rect 572858 480 573830 536
rect 574054 480 575026 536
rect 575250 480 576222 536
rect 576446 480 577326 536
rect 577550 480 578522 536
rect 578746 480 579718 536
rect 579942 480 580914 536
rect 581138 480 582110 536
rect 582334 480 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583520 701793
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 2143 583520 6260
<< metal4 >>
rect -8576 -7504 -7976 711440
rect -7636 -6564 -7036 710500
rect -6696 -5624 -6096 709560
rect -5756 -4684 -5156 708620
rect -4816 -3744 -4216 707680
rect -3876 -2804 -3276 706740
rect -2936 -1864 -2336 705800
rect -1996 -924 -1396 704860
rect 1804 -1864 2404 705800
rect 5404 -3744 6004 707680
rect 9004 -5624 9604 709560
rect 12604 -7504 13204 711440
rect 19804 -1864 20404 705800
rect 23404 -3744 24004 707680
rect 27004 -5624 27604 709560
rect 30604 -7504 31204 711440
rect 37804 666052 38404 705800
rect 41404 666100 42004 707680
rect 45004 666100 45604 709560
rect 48604 666100 49204 711440
rect 55804 666052 56404 705800
rect 59404 666100 60004 707680
rect 63004 666100 63604 709560
rect 66604 666100 67204 711440
rect 73804 666052 74404 705800
rect 77404 666100 78004 707680
rect 81004 666100 81604 709560
rect 84604 666100 85204 711440
rect 91804 666052 92404 705800
rect 95404 666100 96004 707680
rect 99004 666100 99604 709560
rect 102604 666100 103204 711440
rect 109804 666052 110404 705800
rect 113404 666100 114004 707680
rect 117004 666100 117604 709560
rect 120604 666100 121204 711440
rect 127804 666052 128404 705800
rect 131404 666100 132004 707680
rect 135004 666100 135604 709560
rect 138604 666100 139204 711440
rect 145804 666052 146404 705800
rect 149404 666100 150004 707680
rect 153004 666100 153604 709560
rect 156604 666100 157204 711440
rect 163804 666052 164404 705800
rect 167404 666100 168004 707680
rect 171004 666100 171604 709560
rect 174604 666100 175204 711440
rect 181804 666052 182404 705800
rect 185404 666100 186004 707680
rect 189004 666100 189604 709560
rect 192604 666100 193204 711440
rect 199804 666052 200404 705800
rect 203404 666100 204004 707680
rect 207004 666100 207604 709560
rect 210604 666100 211204 711440
rect 217804 666052 218404 705800
rect 221404 666100 222004 707680
rect 225004 666100 225604 709560
rect 228604 666100 229204 711440
rect 235804 666052 236404 705800
rect 239404 666100 240004 707680
rect 243004 666100 243604 709560
rect 246604 666100 247204 711440
rect 253804 666052 254404 705800
rect 257404 666100 258004 707680
rect 37804 495716 38404 518048
rect 41404 495764 42004 518000
rect 45004 495764 45604 518000
rect 48604 495764 49204 518000
rect 55804 495716 56404 518048
rect 59404 495764 60004 518000
rect 63004 495764 63604 518000
rect 66604 495764 67204 518000
rect 73804 495716 74404 518048
rect 77404 495764 78004 518000
rect 81004 495764 81604 518000
rect 84604 495764 85204 518000
rect 91804 495716 92404 518048
rect 95404 495764 96004 518000
rect 99004 495764 99604 518000
rect 102604 495764 103204 518000
rect 109804 495716 110404 518048
rect 113404 495764 114004 518000
rect 117004 495764 117604 518000
rect 120604 495764 121204 518000
rect 127804 495716 128404 518048
rect 131404 495764 132004 518000
rect 135004 495764 135604 518000
rect 138604 495764 139204 518000
rect 145804 495716 146404 518048
rect 149404 495764 150004 518000
rect 153004 495764 153604 518000
rect 156604 495764 157204 518000
rect 163804 495716 164404 518048
rect 167404 495764 168004 518000
rect 171004 495764 171604 518000
rect 174604 495764 175204 518000
rect 37804 325260 38404 358048
rect 41404 325308 42004 358000
rect 45004 325308 45604 358000
rect 48604 325308 49204 358000
rect 55804 325260 56404 358048
rect 59404 325308 60004 358000
rect 63004 325308 63604 358000
rect 66604 325308 67204 358000
rect 73804 325260 74404 358048
rect 77404 325308 78004 358000
rect 81004 325308 81604 358000
rect 84604 325308 85204 358000
rect 91804 325260 92404 358048
rect 95404 325308 96004 358000
rect 99004 325308 99604 358000
rect 102604 325308 103204 358000
rect 109804 325260 110404 358048
rect 113404 325308 114004 358000
rect 117004 325308 117604 358000
rect 120604 325308 121204 358000
rect 127804 325260 128404 358048
rect 131404 325308 132004 358000
rect 135004 325308 135604 358000
rect 138604 325308 139204 358000
rect 145804 325260 146404 358048
rect 149404 325308 150004 358000
rect 153004 325308 153604 358000
rect 156604 325308 157204 358000
rect 163804 325260 164404 358048
rect 167404 325308 168004 358000
rect 171004 325308 171604 358000
rect 174604 325308 175204 358000
rect 37804 221452 38404 238048
rect 41404 221500 42004 238000
rect 45004 221500 45604 238000
rect 48604 221500 49204 238000
rect 55804 221452 56404 238048
rect 59404 221500 60004 238000
rect 63004 221500 63604 238000
rect 66604 221500 67204 238000
rect 73804 221452 74404 238048
rect 77404 221500 78004 238000
rect 81004 221500 81604 238000
rect 84604 221500 85204 238000
rect 91804 221452 92404 238048
rect 95404 221500 96004 238000
rect 99004 221500 99604 238000
rect 102604 221500 103204 238000
rect 109804 221452 110404 238048
rect 113404 221500 114004 238000
rect 117004 221500 117604 238000
rect 120604 221500 121204 238000
rect 127804 221452 128404 238048
rect 131404 221500 132004 238000
rect 135004 221500 135604 238000
rect 37804 111244 38404 138048
rect 41404 111292 42004 138000
rect 45004 111292 45604 138000
rect 48604 111292 49204 138000
rect 55804 111244 56404 138048
rect 59404 111292 60004 138000
rect 63004 111292 63604 138000
rect 66604 111292 67204 138000
rect 73804 111244 74404 138048
rect 77404 111292 78004 138000
rect 81004 111292 81604 138000
rect 84604 111292 85204 138000
rect 91804 111244 92404 138048
rect 95404 111292 96004 138000
rect 99004 111292 99604 138000
rect 102604 111292 103204 138000
rect 109804 111244 110404 138048
rect 113404 111292 114004 138000
rect 117004 111292 117604 138000
rect 120604 111292 121204 138000
rect 127804 111244 128404 138048
rect 131404 111292 132004 138000
rect 37804 -1864 38404 18048
rect 41404 -3744 42004 18000
rect 45004 -5624 45604 18000
rect 48604 -7504 49204 18000
rect 55804 -1864 56404 18048
rect 59404 -3744 60004 18000
rect 63004 -5624 63604 18000
rect 66604 -7504 67204 18000
rect 73804 -1864 74404 18048
rect 77404 -3744 78004 18000
rect 81004 -5624 81604 18000
rect 84604 -7504 85204 18000
rect 91804 -1864 92404 18048
rect 95404 -3744 96004 18000
rect 99004 -5624 99604 18000
rect 102604 -7504 103204 18000
rect 109804 -1864 110404 18048
rect 113404 -3744 114004 18000
rect 117004 -5624 117604 18000
rect 120604 -7504 121204 18000
rect 127804 -1864 128404 18048
rect 131404 -3744 132004 18000
rect 135004 -5624 135604 138000
rect 138604 -7504 139204 238000
rect 145804 -1864 146404 238048
rect 149404 -3744 150004 238000
rect 153004 -5624 153604 238000
rect 156604 -7504 157204 238000
rect 163804 -1864 164404 238048
rect 167404 -3744 168004 238000
rect 171004 -5624 171604 238000
rect 174604 -7504 175204 238000
rect 181804 -1864 182404 518048
rect 185404 -3744 186004 518000
rect 189004 -5624 189604 518000
rect 192604 -7504 193204 518000
rect 199804 -1864 200404 518048
rect 203404 -3744 204004 518000
rect 207004 -5624 207604 518000
rect 210604 -7504 211204 518000
rect 217804 -1864 218404 518048
rect 221404 -3744 222004 518000
rect 225004 -5624 225604 518000
rect 228604 -7504 229204 518000
rect 235804 -1864 236404 518048
rect 239404 -3744 240004 518000
rect 243004 -5624 243604 518000
rect 246604 -7504 247204 518000
rect 253804 -1864 254404 518048
rect 257404 -3744 258004 518000
rect 261004 -5624 261604 709560
rect 264604 -7504 265204 711440
rect 271804 -1864 272404 705800
rect 275404 -3744 276004 707680
rect 279004 -5624 279604 709560
rect 282604 -7504 283204 711440
rect 289804 -1864 290404 705800
rect 293404 -3744 294004 707680
rect 297004 -5624 297604 709560
rect 300604 -7504 301204 711440
rect 307804 -1864 308404 705800
rect 311404 -3744 312004 707680
rect 315004 -5624 315604 709560
rect 318604 -7504 319204 711440
rect 325804 -1864 326404 705800
rect 329404 -3744 330004 707680
rect 333004 -5624 333604 709560
rect 336604 -7504 337204 711440
rect 343804 -1864 344404 705800
rect 347404 -3744 348004 707680
rect 351004 -5624 351604 709560
rect 354604 -7504 355204 711440
rect 361804 -1864 362404 705800
rect 365404 -3744 366004 707680
rect 369004 -5624 369604 709560
rect 372604 -7504 373204 711440
rect 379804 -1864 380404 705800
rect 383404 -3744 384004 707680
rect 387004 -5624 387604 709560
rect 390604 -7504 391204 711440
rect 397804 565820 398404 705800
rect 401404 565868 402004 707680
rect 405004 565868 405604 709560
rect 408604 565868 409204 711440
rect 415804 565820 416404 705800
rect 419404 565868 420004 707680
rect 423004 565868 423604 709560
rect 426604 565868 427204 711440
rect 433804 565820 434404 705800
rect 437404 565868 438004 707680
rect 441004 565868 441604 709560
rect 444604 565868 445204 711440
rect 451804 565820 452404 705800
rect 455404 565868 456004 707680
rect 459004 565868 459604 709560
rect 462604 565868 463204 711440
rect 469804 565820 470404 705800
rect 473404 565868 474004 707680
rect 477004 565868 477604 709560
rect 480604 565868 481204 711440
rect 487804 565820 488404 705800
rect 491404 565868 492004 707680
rect 495004 565868 495604 709560
rect 397804 425812 398404 518048
rect 401404 425860 402004 518000
rect 405004 425860 405604 518000
rect 408604 425860 409204 518000
rect 415804 425812 416404 518048
rect 419404 425860 420004 518000
rect 423004 425860 423604 518000
rect 426604 425860 427204 518000
rect 433804 425812 434404 518048
rect 437404 425860 438004 518000
rect 441004 425860 441604 518000
rect 444604 425860 445204 518000
rect 451804 425812 452404 518048
rect 455404 425860 456004 518000
rect 459004 425860 459604 518000
rect 462604 425860 463204 518000
rect 469804 425812 470404 518048
rect 473404 425860 474004 518000
rect 477004 425860 477604 518000
rect 480604 425860 481204 518000
rect 487804 425812 488404 518048
rect 491404 425860 492004 518000
rect 495004 425860 495604 518000
rect 397804 311388 398404 358048
rect 401404 311436 402004 358000
rect 405004 311436 405604 358000
rect 408604 311436 409204 358000
rect 415804 311388 416404 358048
rect 419404 311436 420004 358000
rect 423004 311436 423604 358000
rect 426604 311436 427204 358000
rect 433804 311388 434404 358048
rect 437404 311436 438004 358000
rect 441004 311436 441604 358000
rect 444604 311436 445204 358000
rect 451804 311388 452404 358048
rect 455404 311436 456004 358000
rect 459004 311436 459604 358000
rect 462604 311436 463204 358000
rect 469804 311388 470404 358048
rect 473404 311436 474004 358000
rect 477004 311436 477604 358000
rect 480604 311436 481204 358000
rect 487804 311388 488404 358048
rect 491404 311436 492004 358000
rect 495004 311436 495604 358000
rect 498604 311436 499204 711440
rect 505804 311388 506404 705800
rect 509404 311436 510004 707680
rect 513004 311436 513604 709560
rect 516604 311436 517204 711440
rect 523804 311388 524404 705800
rect 527404 311436 528004 707680
rect 531004 311436 531604 709560
rect 534604 311436 535204 711440
rect 541804 311388 542404 705800
rect 545404 311436 546004 707680
rect 549004 311436 549604 709560
rect 552604 311436 553204 711440
rect 559804 311388 560404 705800
rect 397804 208940 398404 238048
rect 401404 208988 402004 238000
rect 405004 208988 405604 238000
rect 408604 208988 409204 238000
rect 415804 208940 416404 238048
rect 419404 208988 420004 238000
rect 423004 208988 423604 238000
rect 426604 208988 427204 238000
rect 433804 208940 434404 238048
rect 437404 208988 438004 238000
rect 441004 208988 441604 238000
rect 444604 208988 445204 238000
rect 451804 208940 452404 238048
rect 455404 208988 456004 238000
rect 459004 208988 459604 238000
rect 462604 208988 463204 238000
rect 469804 208940 470404 238048
rect 473404 208988 474004 238000
rect 477004 208988 477604 238000
rect 480604 208988 481204 238000
rect 487804 208940 488404 238048
rect 491404 208988 492004 238000
rect 495004 208988 495604 238000
rect 498604 208988 499204 238000
rect 505804 208940 506404 238048
rect 509404 208988 510004 238000
rect 513004 208988 513604 238000
rect 516604 208988 517204 238000
rect 523804 208940 524404 238048
rect 527404 208988 528004 238000
rect 531004 208988 531604 238000
rect 534604 208988 535204 238000
rect 541804 208940 542404 238048
rect 545404 208988 546004 238000
rect 549004 208988 549604 238000
rect 552604 208988 553204 238000
rect 559804 208940 560404 238048
rect 563404 208988 564004 707680
rect 397804 -1864 398404 138048
rect 401404 -3744 402004 138000
rect 405004 -5624 405604 138000
rect 408604 -7504 409204 138000
rect 415804 -1864 416404 138048
rect 419404 -3744 420004 138000
rect 423004 -5624 423604 138000
rect 426604 -7504 427204 138000
rect 433804 -1864 434404 138048
rect 437404 -3744 438004 138000
rect 441004 -5624 441604 138000
rect 444604 -7504 445204 138000
rect 451804 -1864 452404 138048
rect 455404 -3744 456004 138000
rect 459004 -5624 459604 138000
rect 462604 -7504 463204 138000
rect 469804 -1864 470404 138048
rect 473404 -3744 474004 138000
rect 477004 -5624 477604 138000
rect 480604 -7504 481204 138000
rect 487804 -1864 488404 138048
rect 491404 -3744 492004 138000
rect 495004 -5624 495604 138000
rect 498604 -7504 499204 138000
rect 505804 -1864 506404 138048
rect 509404 -3744 510004 138000
rect 513004 -5624 513604 138000
rect 516604 -7504 517204 138000
rect 523804 -1864 524404 138048
rect 527404 -3744 528004 138000
rect 531004 -5624 531604 138000
rect 534604 -7504 535204 138000
rect 541804 -1864 542404 138048
rect 545404 -3744 546004 138000
rect 549004 -5624 549604 138000
rect 552604 -7504 553204 138000
rect 559804 -1864 560404 138048
rect 563404 -3744 564004 138000
rect 567004 -5624 567604 709560
rect 570604 -7504 571204 711440
rect 577804 -1864 578404 705800
rect 581404 -3744 582004 707680
rect 585320 -924 585920 704860
rect 586260 -1864 586860 705800
rect 587200 -2804 587800 706740
rect 588140 -3744 588740 707680
rect 589080 -4684 589680 708620
rect 590020 -5624 590620 709560
rect 590960 -6564 591560 710500
rect 591900 -7504 592500 711440
<< obsm4 >>
rect 34283 665972 37724 700365
rect 38484 666020 41324 700365
rect 42084 666020 44924 700365
rect 45684 666020 48524 700365
rect 49284 666020 55724 700365
rect 38484 665972 55724 666020
rect 56484 666020 59324 700365
rect 60084 666020 62924 700365
rect 63684 666020 66524 700365
rect 67284 666020 73724 700365
rect 56484 665972 73724 666020
rect 74484 666020 77324 700365
rect 78084 666020 80924 700365
rect 81684 666020 84524 700365
rect 85284 666020 91724 700365
rect 74484 665972 91724 666020
rect 92484 666020 95324 700365
rect 96084 666020 98924 700365
rect 99684 666020 102524 700365
rect 103284 666020 109724 700365
rect 92484 665972 109724 666020
rect 110484 666020 113324 700365
rect 114084 666020 116924 700365
rect 117684 666020 120524 700365
rect 121284 666020 127724 700365
rect 110484 665972 127724 666020
rect 128484 666020 131324 700365
rect 132084 666020 134924 700365
rect 135684 666020 138524 700365
rect 139284 666020 145724 700365
rect 128484 665972 145724 666020
rect 146484 666020 149324 700365
rect 150084 666020 152924 700365
rect 153684 666020 156524 700365
rect 157284 666020 163724 700365
rect 146484 665972 163724 666020
rect 164484 666020 167324 700365
rect 168084 666020 170924 700365
rect 171684 666020 174524 700365
rect 175284 666020 181724 700365
rect 164484 665972 181724 666020
rect 182484 666020 185324 700365
rect 186084 666020 188924 700365
rect 189684 666020 192524 700365
rect 193284 666020 199724 700365
rect 182484 665972 199724 666020
rect 200484 666020 203324 700365
rect 204084 666020 206924 700365
rect 207684 666020 210524 700365
rect 211284 666020 217724 700365
rect 200484 665972 217724 666020
rect 218484 666020 221324 700365
rect 222084 666020 224924 700365
rect 225684 666020 228524 700365
rect 229284 666020 235724 700365
rect 218484 665972 235724 666020
rect 236484 666020 239324 700365
rect 240084 666020 242924 700365
rect 243684 666020 246524 700365
rect 247284 666020 253724 700365
rect 236484 665972 253724 666020
rect 254484 666020 257324 700365
rect 258084 666020 260924 700365
rect 254484 665972 260924 666020
rect 34283 518128 260924 665972
rect 34283 495636 37724 518128
rect 38484 518080 55724 518128
rect 38484 495684 41324 518080
rect 42084 495684 44924 518080
rect 45684 495684 48524 518080
rect 49284 495684 55724 518080
rect 56484 518080 73724 518128
rect 38484 495636 55724 495684
rect 56484 495684 59324 518080
rect 60084 495684 62924 518080
rect 63684 495684 66524 518080
rect 67284 495684 73724 518080
rect 74484 518080 91724 518128
rect 56484 495636 73724 495684
rect 74484 495684 77324 518080
rect 78084 495684 80924 518080
rect 81684 495684 84524 518080
rect 85284 495684 91724 518080
rect 92484 518080 109724 518128
rect 74484 495636 91724 495684
rect 92484 495684 95324 518080
rect 96084 495684 98924 518080
rect 99684 495684 102524 518080
rect 103284 495684 109724 518080
rect 110484 518080 127724 518128
rect 92484 495636 109724 495684
rect 110484 495684 113324 518080
rect 114084 495684 116924 518080
rect 117684 495684 120524 518080
rect 121284 495684 127724 518080
rect 128484 518080 145724 518128
rect 110484 495636 127724 495684
rect 128484 495684 131324 518080
rect 132084 495684 134924 518080
rect 135684 495684 138524 518080
rect 139284 495684 145724 518080
rect 146484 518080 163724 518128
rect 128484 495636 145724 495684
rect 146484 495684 149324 518080
rect 150084 495684 152924 518080
rect 153684 495684 156524 518080
rect 157284 495684 163724 518080
rect 164484 518080 181724 518128
rect 146484 495636 163724 495684
rect 164484 495684 167324 518080
rect 168084 495684 170924 518080
rect 171684 495684 174524 518080
rect 175284 495684 181724 518080
rect 182484 518080 199724 518128
rect 164484 495636 181724 495684
rect 34283 358128 181724 495636
rect 34283 325180 37724 358128
rect 38484 358080 55724 358128
rect 38484 325228 41324 358080
rect 42084 325228 44924 358080
rect 45684 325228 48524 358080
rect 49284 325228 55724 358080
rect 56484 358080 73724 358128
rect 38484 325180 55724 325228
rect 56484 325228 59324 358080
rect 60084 325228 62924 358080
rect 63684 325228 66524 358080
rect 67284 325228 73724 358080
rect 74484 358080 91724 358128
rect 56484 325180 73724 325228
rect 74484 325228 77324 358080
rect 78084 325228 80924 358080
rect 81684 325228 84524 358080
rect 85284 325228 91724 358080
rect 92484 358080 109724 358128
rect 74484 325180 91724 325228
rect 92484 325228 95324 358080
rect 96084 325228 98924 358080
rect 99684 325228 102524 358080
rect 103284 325228 109724 358080
rect 110484 358080 127724 358128
rect 92484 325180 109724 325228
rect 110484 325228 113324 358080
rect 114084 325228 116924 358080
rect 117684 325228 120524 358080
rect 121284 325228 127724 358080
rect 128484 358080 145724 358128
rect 110484 325180 127724 325228
rect 128484 325228 131324 358080
rect 132084 325228 134924 358080
rect 135684 325228 138524 358080
rect 139284 325228 145724 358080
rect 146484 358080 163724 358128
rect 128484 325180 145724 325228
rect 146484 325228 149324 358080
rect 150084 325228 152924 358080
rect 153684 325228 156524 358080
rect 157284 325228 163724 358080
rect 164484 358080 181724 358128
rect 146484 325180 163724 325228
rect 164484 325228 167324 358080
rect 168084 325228 170924 358080
rect 171684 325228 174524 358080
rect 175284 325228 181724 358080
rect 164484 325180 181724 325228
rect 34283 238128 181724 325180
rect 34283 221372 37724 238128
rect 38484 238080 55724 238128
rect 38484 221420 41324 238080
rect 42084 221420 44924 238080
rect 45684 221420 48524 238080
rect 49284 221420 55724 238080
rect 56484 238080 73724 238128
rect 38484 221372 55724 221420
rect 56484 221420 59324 238080
rect 60084 221420 62924 238080
rect 63684 221420 66524 238080
rect 67284 221420 73724 238080
rect 74484 238080 91724 238128
rect 56484 221372 73724 221420
rect 74484 221420 77324 238080
rect 78084 221420 80924 238080
rect 81684 221420 84524 238080
rect 85284 221420 91724 238080
rect 92484 238080 109724 238128
rect 74484 221372 91724 221420
rect 92484 221420 95324 238080
rect 96084 221420 98924 238080
rect 99684 221420 102524 238080
rect 103284 221420 109724 238080
rect 110484 238080 127724 238128
rect 92484 221372 109724 221420
rect 110484 221420 113324 238080
rect 114084 221420 116924 238080
rect 117684 221420 120524 238080
rect 121284 221420 127724 238080
rect 128484 238080 145724 238128
rect 110484 221372 127724 221420
rect 128484 221420 131324 238080
rect 132084 221420 134924 238080
rect 135684 221420 138524 238080
rect 128484 221372 138524 221420
rect 34283 138128 138524 221372
rect 34283 111164 37724 138128
rect 38484 138080 55724 138128
rect 38484 111212 41324 138080
rect 42084 111212 44924 138080
rect 45684 111212 48524 138080
rect 49284 111212 55724 138080
rect 56484 138080 73724 138128
rect 38484 111164 55724 111212
rect 56484 111212 59324 138080
rect 60084 111212 62924 138080
rect 63684 111212 66524 138080
rect 67284 111212 73724 138080
rect 74484 138080 91724 138128
rect 56484 111164 73724 111212
rect 74484 111212 77324 138080
rect 78084 111212 80924 138080
rect 81684 111212 84524 138080
rect 85284 111212 91724 138080
rect 92484 138080 109724 138128
rect 74484 111164 91724 111212
rect 92484 111212 95324 138080
rect 96084 111212 98924 138080
rect 99684 111212 102524 138080
rect 103284 111212 109724 138080
rect 110484 138080 127724 138128
rect 92484 111164 109724 111212
rect 110484 111212 113324 138080
rect 114084 111212 116924 138080
rect 117684 111212 120524 138080
rect 121284 111212 127724 138080
rect 128484 138080 138524 138128
rect 110484 111164 127724 111212
rect 128484 111212 131324 138080
rect 132084 111212 134924 138080
rect 128484 111164 134924 111212
rect 34283 18128 134924 111164
rect 34283 3027 37724 18128
rect 38484 18080 55724 18128
rect 38484 3027 41324 18080
rect 42084 3027 44924 18080
rect 45684 3027 48524 18080
rect 49284 3027 55724 18080
rect 56484 18080 73724 18128
rect 56484 3027 59324 18080
rect 60084 3027 62924 18080
rect 63684 3027 66524 18080
rect 67284 3027 73724 18080
rect 74484 18080 91724 18128
rect 74484 3027 77324 18080
rect 78084 3027 80924 18080
rect 81684 3027 84524 18080
rect 85284 3027 91724 18080
rect 92484 18080 109724 18128
rect 92484 3027 95324 18080
rect 96084 3027 98924 18080
rect 99684 3027 102524 18080
rect 103284 3027 109724 18080
rect 110484 18080 127724 18128
rect 110484 3027 113324 18080
rect 114084 3027 116924 18080
rect 117684 3027 120524 18080
rect 121284 3027 127724 18080
rect 128484 18080 134924 18128
rect 128484 3027 131324 18080
rect 132084 3027 134924 18080
rect 135684 3027 138524 138080
rect 139284 3027 145724 238080
rect 146484 238080 163724 238128
rect 146484 3027 149324 238080
rect 150084 3027 152924 238080
rect 153684 3027 156524 238080
rect 157284 3027 163724 238080
rect 164484 238080 181724 238128
rect 164484 3027 167324 238080
rect 168084 3027 170924 238080
rect 171684 3027 174524 238080
rect 175284 3027 181724 238080
rect 182484 3027 185324 518080
rect 186084 3027 188924 518080
rect 189684 3027 192524 518080
rect 193284 3027 199724 518080
rect 200484 518080 217724 518128
rect 200484 3027 203324 518080
rect 204084 3027 206924 518080
rect 207684 3027 210524 518080
rect 211284 3027 217724 518080
rect 218484 518080 235724 518128
rect 218484 3027 221324 518080
rect 222084 3027 224924 518080
rect 225684 3027 228524 518080
rect 229284 3027 235724 518080
rect 236484 518080 253724 518128
rect 236484 3027 239324 518080
rect 240084 3027 242924 518080
rect 243684 3027 246524 518080
rect 247284 3027 253724 518080
rect 254484 518080 260924 518128
rect 254484 3027 257324 518080
rect 258084 3027 260924 518080
rect 261684 3027 264524 700365
rect 265284 3027 271724 700365
rect 272484 3027 275324 700365
rect 276084 3027 278924 700365
rect 279684 3027 282524 700365
rect 283284 3027 289724 700365
rect 290484 3027 293324 700365
rect 294084 3027 296924 700365
rect 297684 3027 300524 700365
rect 301284 3027 307724 700365
rect 308484 3027 311324 700365
rect 312084 3027 314924 700365
rect 315684 3027 318524 700365
rect 319284 3027 325724 700365
rect 326484 3027 329324 700365
rect 330084 3027 332924 700365
rect 333684 3027 336524 700365
rect 337284 3027 343724 700365
rect 344484 3027 347324 700365
rect 348084 3027 350924 700365
rect 351684 3027 354524 700365
rect 355284 3027 361724 700365
rect 362484 3027 365324 700365
rect 366084 3027 368924 700365
rect 369684 3027 372524 700365
rect 373284 3027 379724 700365
rect 380484 3027 383324 700365
rect 384084 3027 386924 700365
rect 387684 3027 390524 700365
rect 391284 565740 397724 700365
rect 398484 565788 401324 700365
rect 402084 565788 404924 700365
rect 405684 565788 408524 700365
rect 409284 565788 415724 700365
rect 398484 565740 415724 565788
rect 416484 565788 419324 700365
rect 420084 565788 422924 700365
rect 423684 565788 426524 700365
rect 427284 565788 433724 700365
rect 416484 565740 433724 565788
rect 434484 565788 437324 700365
rect 438084 565788 440924 700365
rect 441684 565788 444524 700365
rect 445284 565788 451724 700365
rect 434484 565740 451724 565788
rect 452484 565788 455324 700365
rect 456084 565788 458924 700365
rect 459684 565788 462524 700365
rect 463284 565788 469724 700365
rect 452484 565740 469724 565788
rect 470484 565788 473324 700365
rect 474084 565788 476924 700365
rect 477684 565788 480524 700365
rect 481284 565788 487724 700365
rect 470484 565740 487724 565788
rect 488484 565788 491324 700365
rect 492084 565788 494924 700365
rect 495684 565788 498524 700365
rect 488484 565740 498524 565788
rect 391284 518128 498524 565740
rect 391284 425732 397724 518128
rect 398484 518080 415724 518128
rect 398484 425780 401324 518080
rect 402084 425780 404924 518080
rect 405684 425780 408524 518080
rect 409284 425780 415724 518080
rect 416484 518080 433724 518128
rect 398484 425732 415724 425780
rect 416484 425780 419324 518080
rect 420084 425780 422924 518080
rect 423684 425780 426524 518080
rect 427284 425780 433724 518080
rect 434484 518080 451724 518128
rect 416484 425732 433724 425780
rect 434484 425780 437324 518080
rect 438084 425780 440924 518080
rect 441684 425780 444524 518080
rect 445284 425780 451724 518080
rect 452484 518080 469724 518128
rect 434484 425732 451724 425780
rect 452484 425780 455324 518080
rect 456084 425780 458924 518080
rect 459684 425780 462524 518080
rect 463284 425780 469724 518080
rect 470484 518080 487724 518128
rect 452484 425732 469724 425780
rect 470484 425780 473324 518080
rect 474084 425780 476924 518080
rect 477684 425780 480524 518080
rect 481284 425780 487724 518080
rect 488484 518080 498524 518128
rect 470484 425732 487724 425780
rect 488484 425780 491324 518080
rect 492084 425780 494924 518080
rect 495684 425780 498524 518080
rect 488484 425732 498524 425780
rect 391284 358128 498524 425732
rect 391284 311308 397724 358128
rect 398484 358080 415724 358128
rect 398484 311356 401324 358080
rect 402084 311356 404924 358080
rect 405684 311356 408524 358080
rect 409284 311356 415724 358080
rect 416484 358080 433724 358128
rect 398484 311308 415724 311356
rect 416484 311356 419324 358080
rect 420084 311356 422924 358080
rect 423684 311356 426524 358080
rect 427284 311356 433724 358080
rect 434484 358080 451724 358128
rect 416484 311308 433724 311356
rect 434484 311356 437324 358080
rect 438084 311356 440924 358080
rect 441684 311356 444524 358080
rect 445284 311356 451724 358080
rect 452484 358080 469724 358128
rect 434484 311308 451724 311356
rect 452484 311356 455324 358080
rect 456084 311356 458924 358080
rect 459684 311356 462524 358080
rect 463284 311356 469724 358080
rect 470484 358080 487724 358128
rect 452484 311308 469724 311356
rect 470484 311356 473324 358080
rect 474084 311356 476924 358080
rect 477684 311356 480524 358080
rect 481284 311356 487724 358080
rect 488484 358080 498524 358128
rect 470484 311308 487724 311356
rect 488484 311356 491324 358080
rect 492084 311356 494924 358080
rect 495684 311356 498524 358080
rect 499284 311356 505724 700365
rect 488484 311308 505724 311356
rect 506484 311356 509324 700365
rect 510084 311356 512924 700365
rect 513684 311356 516524 700365
rect 517284 311356 523724 700365
rect 506484 311308 523724 311356
rect 524484 311356 527324 700365
rect 528084 311356 530924 700365
rect 531684 311356 534524 700365
rect 535284 311356 541724 700365
rect 524484 311308 541724 311356
rect 542484 311356 545324 700365
rect 546084 311356 548924 700365
rect 549684 311356 552524 700365
rect 553284 311356 559724 700365
rect 542484 311308 559724 311356
rect 560484 311308 563324 700365
rect 391284 238128 563324 311308
rect 391284 208860 397724 238128
rect 398484 238080 415724 238128
rect 398484 208908 401324 238080
rect 402084 208908 404924 238080
rect 405684 208908 408524 238080
rect 409284 208908 415724 238080
rect 416484 238080 433724 238128
rect 398484 208860 415724 208908
rect 416484 208908 419324 238080
rect 420084 208908 422924 238080
rect 423684 208908 426524 238080
rect 427284 208908 433724 238080
rect 434484 238080 451724 238128
rect 416484 208860 433724 208908
rect 434484 208908 437324 238080
rect 438084 208908 440924 238080
rect 441684 208908 444524 238080
rect 445284 208908 451724 238080
rect 452484 238080 469724 238128
rect 434484 208860 451724 208908
rect 452484 208908 455324 238080
rect 456084 208908 458924 238080
rect 459684 208908 462524 238080
rect 463284 208908 469724 238080
rect 470484 238080 487724 238128
rect 452484 208860 469724 208908
rect 470484 208908 473324 238080
rect 474084 208908 476924 238080
rect 477684 208908 480524 238080
rect 481284 208908 487724 238080
rect 488484 238080 505724 238128
rect 470484 208860 487724 208908
rect 488484 208908 491324 238080
rect 492084 208908 494924 238080
rect 495684 208908 498524 238080
rect 499284 208908 505724 238080
rect 506484 238080 523724 238128
rect 488484 208860 505724 208908
rect 506484 208908 509324 238080
rect 510084 208908 512924 238080
rect 513684 208908 516524 238080
rect 517284 208908 523724 238080
rect 524484 238080 541724 238128
rect 506484 208860 523724 208908
rect 524484 208908 527324 238080
rect 528084 208908 530924 238080
rect 531684 208908 534524 238080
rect 535284 208908 541724 238080
rect 542484 238080 559724 238128
rect 524484 208860 541724 208908
rect 542484 208908 545324 238080
rect 546084 208908 548924 238080
rect 549684 208908 552524 238080
rect 553284 208908 559724 238080
rect 542484 208860 559724 208908
rect 560484 208908 563324 238128
rect 564084 208908 564376 700365
rect 560484 208860 564376 208908
rect 391284 138128 564376 208860
rect 391284 3027 397724 138128
rect 398484 138080 415724 138128
rect 398484 3027 401324 138080
rect 402084 3027 404924 138080
rect 405684 3027 408524 138080
rect 409284 3027 415724 138080
rect 416484 138080 433724 138128
rect 416484 3027 419324 138080
rect 420084 3027 422924 138080
rect 423684 3027 426524 138080
rect 427284 3027 433724 138080
rect 434484 138080 451724 138128
rect 434484 3027 437324 138080
rect 438084 3027 440924 138080
rect 441684 3027 444524 138080
rect 445284 3027 451724 138080
rect 452484 138080 469724 138128
rect 452484 3027 455324 138080
rect 456084 3027 458924 138080
rect 459684 3027 462524 138080
rect 463284 3027 469724 138080
rect 470484 138080 487724 138128
rect 470484 3027 473324 138080
rect 474084 3027 476924 138080
rect 477684 3027 480524 138080
rect 481284 3027 487724 138080
rect 488484 138080 505724 138128
rect 488484 3027 491324 138080
rect 492084 3027 494924 138080
rect 495684 3027 498524 138080
rect 499284 3027 505724 138080
rect 506484 138080 523724 138128
rect 506484 3027 509324 138080
rect 510084 3027 512924 138080
rect 513684 3027 516524 138080
rect 517284 3027 523724 138080
rect 524484 138080 541724 138128
rect 524484 3027 527324 138080
rect 528084 3027 530924 138080
rect 531684 3027 534524 138080
rect 535284 3027 541724 138080
rect 542484 138080 559724 138128
rect 542484 3027 545324 138080
rect 546084 3027 548924 138080
rect 549684 3027 552524 138080
rect 553284 3027 559724 138080
rect 560484 138080 564376 138128
rect 560484 3027 563324 138080
rect 564084 3027 564376 138080
<< metal5 >>
rect -8576 710840 592500 711440
rect -7636 709900 591560 710500
rect -6696 708960 590620 709560
rect -5756 708020 589680 708620
rect -4816 707080 588740 707680
rect -3876 706140 587800 706740
rect -2936 705200 586860 705800
rect -1996 704260 585920 704860
rect -8576 697676 592500 698276
rect -6696 694076 590620 694676
rect -4816 690476 588740 691076
rect -2936 686828 586860 687428
rect -8576 679676 592500 680276
rect -6696 676076 590620 676676
rect -4816 672476 588740 673076
rect -2936 668828 586860 669428
rect -8576 661676 592500 662276
rect -6696 658076 590620 658676
rect -4816 654476 588740 655076
rect -2936 650828 586860 651428
rect -8576 643676 592500 644276
rect -6696 640076 590620 640676
rect -4816 636476 588740 637076
rect -2936 632828 586860 633428
rect -8576 625676 592500 626276
rect -6696 622076 590620 622676
rect -4816 618476 588740 619076
rect -2936 614828 586860 615428
rect -8576 607676 592500 608276
rect -6696 604076 590620 604676
rect -4816 600476 588740 601076
rect -2936 596828 586860 597428
rect -8576 589676 592500 590276
rect -6696 586076 590620 586676
rect -4816 582476 588740 583076
rect -2936 578828 586860 579428
rect -8576 571676 592500 572276
rect -6696 568076 590620 568676
rect -4816 564476 588740 565076
rect -2936 560828 586860 561428
rect -8576 553676 592500 554276
rect -6696 550076 590620 550676
rect -4816 546476 588740 547076
rect -2936 542828 586860 543428
rect -8576 535676 592500 536276
rect -6696 532076 590620 532676
rect -4816 528476 588740 529076
rect -2936 524828 586860 525428
rect -8576 517676 592500 518276
rect -6696 514076 590620 514676
rect -4816 510476 588740 511076
rect -2936 506828 586860 507428
rect -8576 499676 592500 500276
rect -6696 496076 590620 496676
rect -4816 492476 588740 493076
rect -2936 488828 586860 489428
rect -8576 481676 592500 482276
rect -6696 478076 590620 478676
rect -4816 474476 588740 475076
rect -2936 470828 586860 471428
rect -8576 463676 592500 464276
rect -6696 460076 590620 460676
rect -4816 456476 588740 457076
rect -2936 452828 586860 453428
rect -8576 445676 592500 446276
rect -6696 442076 590620 442676
rect -4816 438476 588740 439076
rect -2936 434828 586860 435428
rect -8576 427676 592500 428276
rect -6696 424076 590620 424676
rect -4816 420476 588740 421076
rect -2936 416828 586860 417428
rect -8576 409676 592500 410276
rect -6696 406076 590620 406676
rect -4816 402476 588740 403076
rect -2936 398828 586860 399428
rect -8576 391676 592500 392276
rect -6696 388076 590620 388676
rect -4816 384476 588740 385076
rect -2936 380828 586860 381428
rect -8576 373676 592500 374276
rect -6696 370076 590620 370676
rect -4816 366476 588740 367076
rect -2936 362828 586860 363428
rect -8576 355676 592500 356276
rect -6696 352076 590620 352676
rect -4816 348476 588740 349076
rect -2936 344828 586860 345428
rect -8576 337676 592500 338276
rect -6696 334076 590620 334676
rect -4816 330476 588740 331076
rect -2936 326828 586860 327428
rect -8576 319676 592500 320276
rect -6696 316076 590620 316676
rect -4816 312476 588740 313076
rect -2936 308828 586860 309428
rect -8576 301676 592500 302276
rect -6696 298076 590620 298676
rect -4816 294476 588740 295076
rect -2936 290828 586860 291428
rect -8576 283676 592500 284276
rect -6696 280076 590620 280676
rect -4816 276476 588740 277076
rect -2936 272828 586860 273428
rect -8576 265676 592500 266276
rect -6696 262076 590620 262676
rect -4816 258476 588740 259076
rect -2936 254828 586860 255428
rect -8576 247676 592500 248276
rect -6696 244076 590620 244676
rect -4816 240476 588740 241076
rect -2936 236828 586860 237428
rect -8576 229676 592500 230276
rect -6696 226076 590620 226676
rect -4816 222476 588740 223076
rect -2936 218828 586860 219428
rect -8576 211676 592500 212276
rect -6696 208076 590620 208676
rect -4816 204476 588740 205076
rect -2936 200828 586860 201428
rect -8576 193676 592500 194276
rect -6696 190076 590620 190676
rect -4816 186476 588740 187076
rect -2936 182828 586860 183428
rect -8576 175676 592500 176276
rect -6696 172076 590620 172676
rect -4816 168476 588740 169076
rect -2936 164828 586860 165428
rect -8576 157676 592500 158276
rect -6696 154076 590620 154676
rect -4816 150476 588740 151076
rect -2936 146828 586860 147428
rect -8576 139676 592500 140276
rect -6696 136076 590620 136676
rect -4816 132476 588740 133076
rect -2936 128828 586860 129428
rect -8576 121676 592500 122276
rect -6696 118076 590620 118676
rect -4816 114476 588740 115076
rect -2936 110828 586860 111428
rect -8576 103676 592500 104276
rect -6696 100076 590620 100676
rect -4816 96476 588740 97076
rect -2936 92828 586860 93428
rect -8576 85676 592500 86276
rect -6696 82076 590620 82676
rect -4816 78476 588740 79076
rect -2936 74828 586860 75428
rect -8576 67676 592500 68276
rect -6696 64076 590620 64676
rect -4816 60476 588740 61076
rect -2936 56828 586860 57428
rect -8576 49676 592500 50276
rect -6696 46076 590620 46676
rect -4816 42476 588740 43076
rect -2936 38828 586860 39428
rect -8576 31676 592500 32276
rect -6696 28076 590620 28676
rect -4816 24476 588740 25076
rect -2936 20828 586860 21428
rect -8576 13676 592500 14276
rect -6696 10076 590620 10676
rect -4816 6476 588740 7076
rect -2936 2828 586860 3428
rect -1996 -924 585920 -324
rect -2936 -1864 586860 -1264
rect -3876 -2804 587800 -2204
rect -4816 -3744 588740 -3144
rect -5756 -4684 589680 -4084
rect -6696 -5624 590620 -5024
rect -7636 -6564 591560 -5964
rect -8576 -7504 592500 -6904
<< obsm5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect 0 698596 584000 703940
rect -7636 698276 -7036 698278
rect 590960 698276 591560 698278
rect -7636 697674 -7036 697676
rect 590960 697674 591560 697676
rect 0 694996 584000 697356
rect -5756 694676 -5156 694678
rect 589080 694676 589680 694678
rect -5756 694074 -5156 694076
rect 589080 694074 589680 694076
rect 0 691396 584000 693756
rect -3876 691076 -3276 691078
rect 587200 691076 587800 691078
rect -3876 690474 -3276 690476
rect 587200 690474 587800 690476
rect 0 687748 584000 690156
rect -1996 687428 -1396 687430
rect 585320 687428 585920 687430
rect -1996 686826 -1396 686828
rect 585320 686826 585920 686828
rect 0 680596 584000 686508
rect -8576 680276 -7976 680278
rect 591900 680276 592500 680278
rect -8576 679674 -7976 679676
rect 591900 679674 592500 679676
rect 0 676996 584000 679356
rect -6696 676676 -6096 676678
rect 590020 676676 590620 676678
rect -6696 676074 -6096 676076
rect 590020 676074 590620 676076
rect 0 673396 584000 675756
rect -4816 673076 -4216 673078
rect 588140 673076 588740 673078
rect -4816 672474 -4216 672476
rect 588140 672474 588740 672476
rect 0 669748 584000 672156
rect -2936 669428 -2336 669430
rect 586260 669428 586860 669430
rect -2936 668826 -2336 668828
rect 586260 668826 586860 668828
rect 0 662596 584000 668508
rect -7636 662276 -7036 662278
rect 590960 662276 591560 662278
rect -7636 661674 -7036 661676
rect 590960 661674 591560 661676
rect 0 658996 584000 661356
rect -5756 658676 -5156 658678
rect 589080 658676 589680 658678
rect -5756 658074 -5156 658076
rect 589080 658074 589680 658076
rect 0 655396 584000 657756
rect -3876 655076 -3276 655078
rect 587200 655076 587800 655078
rect -3876 654474 -3276 654476
rect 587200 654474 587800 654476
rect 0 651748 584000 654156
rect -1996 651428 -1396 651430
rect 585320 651428 585920 651430
rect -1996 650826 -1396 650828
rect 585320 650826 585920 650828
rect 0 644596 584000 650508
rect -8576 644276 -7976 644278
rect 591900 644276 592500 644278
rect -8576 643674 -7976 643676
rect 591900 643674 592500 643676
rect 0 640996 584000 643356
rect -6696 640676 -6096 640678
rect 590020 640676 590620 640678
rect -6696 640074 -6096 640076
rect 590020 640074 590620 640076
rect 0 637396 584000 639756
rect -4816 637076 -4216 637078
rect 588140 637076 588740 637078
rect -4816 636474 -4216 636476
rect 588140 636474 588740 636476
rect 0 633748 584000 636156
rect -2936 633428 -2336 633430
rect 586260 633428 586860 633430
rect -2936 632826 -2336 632828
rect 586260 632826 586860 632828
rect 0 626596 584000 632508
rect -7636 626276 -7036 626278
rect 590960 626276 591560 626278
rect -7636 625674 -7036 625676
rect 590960 625674 591560 625676
rect 0 622996 584000 625356
rect -5756 622676 -5156 622678
rect 589080 622676 589680 622678
rect -5756 622074 -5156 622076
rect 589080 622074 589680 622076
rect 0 619396 584000 621756
rect -3876 619076 -3276 619078
rect 587200 619076 587800 619078
rect -3876 618474 -3276 618476
rect 587200 618474 587800 618476
rect 0 615748 584000 618156
rect -1996 615428 -1396 615430
rect 585320 615428 585920 615430
rect -1996 614826 -1396 614828
rect 585320 614826 585920 614828
rect 0 608596 584000 614508
rect -8576 608276 -7976 608278
rect 591900 608276 592500 608278
rect -8576 607674 -7976 607676
rect 591900 607674 592500 607676
rect 0 604996 584000 607356
rect -6696 604676 -6096 604678
rect 590020 604676 590620 604678
rect -6696 604074 -6096 604076
rect 590020 604074 590620 604076
rect 0 601396 584000 603756
rect -4816 601076 -4216 601078
rect 588140 601076 588740 601078
rect -4816 600474 -4216 600476
rect 588140 600474 588740 600476
rect 0 597748 584000 600156
rect -2936 597428 -2336 597430
rect 586260 597428 586860 597430
rect -2936 596826 -2336 596828
rect 586260 596826 586860 596828
rect 0 590596 584000 596508
rect -7636 590276 -7036 590278
rect 590960 590276 591560 590278
rect -7636 589674 -7036 589676
rect 590960 589674 591560 589676
rect 0 586996 584000 589356
rect -5756 586676 -5156 586678
rect 589080 586676 589680 586678
rect -5756 586074 -5156 586076
rect 589080 586074 589680 586076
rect 0 583396 584000 585756
rect -3876 583076 -3276 583078
rect 587200 583076 587800 583078
rect -3876 582474 -3276 582476
rect 587200 582474 587800 582476
rect 0 579748 584000 582156
rect -1996 579428 -1396 579430
rect 585320 579428 585920 579430
rect -1996 578826 -1396 578828
rect 585320 578826 585920 578828
rect 0 572596 584000 578508
rect -8576 572276 -7976 572278
rect 591900 572276 592500 572278
rect -8576 571674 -7976 571676
rect 591900 571674 592500 571676
rect 0 568996 584000 571356
rect -6696 568676 -6096 568678
rect 590020 568676 590620 568678
rect -6696 568074 -6096 568076
rect 590020 568074 590620 568076
rect 0 565396 584000 567756
rect -4816 565076 -4216 565078
rect 588140 565076 588740 565078
rect -4816 564474 -4216 564476
rect 588140 564474 588740 564476
rect 0 561748 584000 564156
rect -2936 561428 -2336 561430
rect 586260 561428 586860 561430
rect -2936 560826 -2336 560828
rect 586260 560826 586860 560828
rect 0 554596 584000 560508
rect -7636 554276 -7036 554278
rect 590960 554276 591560 554278
rect -7636 553674 -7036 553676
rect 590960 553674 591560 553676
rect 0 550996 584000 553356
rect -5756 550676 -5156 550678
rect 589080 550676 589680 550678
rect -5756 550074 -5156 550076
rect 589080 550074 589680 550076
rect 0 547396 584000 549756
rect -3876 547076 -3276 547078
rect 587200 547076 587800 547078
rect -3876 546474 -3276 546476
rect 587200 546474 587800 546476
rect 0 543748 584000 546156
rect -1996 543428 -1396 543430
rect 585320 543428 585920 543430
rect -1996 542826 -1396 542828
rect 585320 542826 585920 542828
rect 0 536596 584000 542508
rect -8576 536276 -7976 536278
rect 591900 536276 592500 536278
rect -8576 535674 -7976 535676
rect 591900 535674 592500 535676
rect 0 532996 584000 535356
rect -6696 532676 -6096 532678
rect 590020 532676 590620 532678
rect -6696 532074 -6096 532076
rect 590020 532074 590620 532076
rect 0 529396 584000 531756
rect -4816 529076 -4216 529078
rect 588140 529076 588740 529078
rect -4816 528474 -4216 528476
rect 588140 528474 588740 528476
rect 0 525748 584000 528156
rect -2936 525428 -2336 525430
rect 586260 525428 586860 525430
rect -2936 524826 -2336 524828
rect 586260 524826 586860 524828
rect 0 518596 584000 524508
rect -7636 518276 -7036 518278
rect 590960 518276 591560 518278
rect -7636 517674 -7036 517676
rect 590960 517674 591560 517676
rect 0 514996 584000 517356
rect -5756 514676 -5156 514678
rect 589080 514676 589680 514678
rect -5756 514074 -5156 514076
rect 589080 514074 589680 514076
rect 0 511396 584000 513756
rect -3876 511076 -3276 511078
rect 587200 511076 587800 511078
rect -3876 510474 -3276 510476
rect 587200 510474 587800 510476
rect 0 507748 584000 510156
rect -1996 507428 -1396 507430
rect 585320 507428 585920 507430
rect -1996 506826 -1396 506828
rect 585320 506826 585920 506828
rect 0 500596 584000 506508
rect -8576 500276 -7976 500278
rect 591900 500276 592500 500278
rect -8576 499674 -7976 499676
rect 591900 499674 592500 499676
rect 0 496996 584000 499356
rect -6696 496676 -6096 496678
rect 590020 496676 590620 496678
rect -6696 496074 -6096 496076
rect 590020 496074 590620 496076
rect 0 493396 584000 495756
rect -4816 493076 -4216 493078
rect 588140 493076 588740 493078
rect -4816 492474 -4216 492476
rect 588140 492474 588740 492476
rect 0 489748 584000 492156
rect -2936 489428 -2336 489430
rect 586260 489428 586860 489430
rect -2936 488826 -2336 488828
rect 586260 488826 586860 488828
rect 0 482596 584000 488508
rect -7636 482276 -7036 482278
rect 590960 482276 591560 482278
rect -7636 481674 -7036 481676
rect 590960 481674 591560 481676
rect 0 478996 584000 481356
rect -5756 478676 -5156 478678
rect 589080 478676 589680 478678
rect -5756 478074 -5156 478076
rect 589080 478074 589680 478076
rect 0 475396 584000 477756
rect -3876 475076 -3276 475078
rect 587200 475076 587800 475078
rect -3876 474474 -3276 474476
rect 587200 474474 587800 474476
rect 0 471748 584000 474156
rect -1996 471428 -1396 471430
rect 585320 471428 585920 471430
rect -1996 470826 -1396 470828
rect 585320 470826 585920 470828
rect 0 464596 584000 470508
rect -8576 464276 -7976 464278
rect 591900 464276 592500 464278
rect -8576 463674 -7976 463676
rect 591900 463674 592500 463676
rect 0 460996 584000 463356
rect -6696 460676 -6096 460678
rect 590020 460676 590620 460678
rect -6696 460074 -6096 460076
rect 590020 460074 590620 460076
rect 0 457396 584000 459756
rect -4816 457076 -4216 457078
rect 588140 457076 588740 457078
rect -4816 456474 -4216 456476
rect 588140 456474 588740 456476
rect 0 453748 584000 456156
rect -2936 453428 -2336 453430
rect 586260 453428 586860 453430
rect -2936 452826 -2336 452828
rect 586260 452826 586860 452828
rect 0 446596 584000 452508
rect -7636 446276 -7036 446278
rect 590960 446276 591560 446278
rect -7636 445674 -7036 445676
rect 590960 445674 591560 445676
rect 0 442996 584000 445356
rect -5756 442676 -5156 442678
rect 589080 442676 589680 442678
rect -5756 442074 -5156 442076
rect 589080 442074 589680 442076
rect 0 439396 584000 441756
rect -3876 439076 -3276 439078
rect 587200 439076 587800 439078
rect -3876 438474 -3276 438476
rect 587200 438474 587800 438476
rect 0 435748 584000 438156
rect -1996 435428 -1396 435430
rect 585320 435428 585920 435430
rect -1996 434826 -1396 434828
rect 585320 434826 585920 434828
rect 0 428596 584000 434508
rect -8576 428276 -7976 428278
rect 591900 428276 592500 428278
rect -8576 427674 -7976 427676
rect 591900 427674 592500 427676
rect 0 424996 584000 427356
rect -6696 424676 -6096 424678
rect 590020 424676 590620 424678
rect -6696 424074 -6096 424076
rect 590020 424074 590620 424076
rect 0 421396 584000 423756
rect -4816 421076 -4216 421078
rect 588140 421076 588740 421078
rect -4816 420474 -4216 420476
rect 588140 420474 588740 420476
rect 0 417748 584000 420156
rect -2936 417428 -2336 417430
rect 586260 417428 586860 417430
rect -2936 416826 -2336 416828
rect 586260 416826 586860 416828
rect 0 410596 584000 416508
rect -7636 410276 -7036 410278
rect 590960 410276 591560 410278
rect -7636 409674 -7036 409676
rect 590960 409674 591560 409676
rect 0 406996 584000 409356
rect -5756 406676 -5156 406678
rect 589080 406676 589680 406678
rect -5756 406074 -5156 406076
rect 589080 406074 589680 406076
rect 0 403396 584000 405756
rect -3876 403076 -3276 403078
rect 587200 403076 587800 403078
rect -3876 402474 -3276 402476
rect 587200 402474 587800 402476
rect 0 399748 584000 402156
rect -1996 399428 -1396 399430
rect 585320 399428 585920 399430
rect -1996 398826 -1396 398828
rect 585320 398826 585920 398828
rect 0 392596 584000 398508
rect -8576 392276 -7976 392278
rect 591900 392276 592500 392278
rect -8576 391674 -7976 391676
rect 591900 391674 592500 391676
rect 0 388996 584000 391356
rect -6696 388676 -6096 388678
rect 590020 388676 590620 388678
rect -6696 388074 -6096 388076
rect 590020 388074 590620 388076
rect 0 385396 584000 387756
rect -4816 385076 -4216 385078
rect 588140 385076 588740 385078
rect -4816 384474 -4216 384476
rect 588140 384474 588740 384476
rect 0 381748 584000 384156
rect -2936 381428 -2336 381430
rect 586260 381428 586860 381430
rect -2936 380826 -2336 380828
rect 586260 380826 586860 380828
rect 0 374596 584000 380508
rect -7636 374276 -7036 374278
rect 590960 374276 591560 374278
rect -7636 373674 -7036 373676
rect 590960 373674 591560 373676
rect 0 370996 584000 373356
rect -5756 370676 -5156 370678
rect 589080 370676 589680 370678
rect -5756 370074 -5156 370076
rect 589080 370074 589680 370076
rect 0 367396 584000 369756
rect -3876 367076 -3276 367078
rect 587200 367076 587800 367078
rect -3876 366474 -3276 366476
rect 587200 366474 587800 366476
rect 0 363748 584000 366156
rect -1996 363428 -1396 363430
rect 585320 363428 585920 363430
rect -1996 362826 -1396 362828
rect 585320 362826 585920 362828
rect 0 356596 584000 362508
rect -8576 356276 -7976 356278
rect 591900 356276 592500 356278
rect -8576 355674 -7976 355676
rect 591900 355674 592500 355676
rect 0 352996 584000 355356
rect -6696 352676 -6096 352678
rect 590020 352676 590620 352678
rect -6696 352074 -6096 352076
rect 590020 352074 590620 352076
rect 0 349396 584000 351756
rect -4816 349076 -4216 349078
rect 588140 349076 588740 349078
rect -4816 348474 -4216 348476
rect 588140 348474 588740 348476
rect 0 345748 584000 348156
rect -2936 345428 -2336 345430
rect 586260 345428 586860 345430
rect -2936 344826 -2336 344828
rect 586260 344826 586860 344828
rect 0 338596 584000 344508
rect -7636 338276 -7036 338278
rect 590960 338276 591560 338278
rect -7636 337674 -7036 337676
rect 590960 337674 591560 337676
rect 0 334996 584000 337356
rect -5756 334676 -5156 334678
rect 589080 334676 589680 334678
rect -5756 334074 -5156 334076
rect 589080 334074 589680 334076
rect 0 331396 584000 333756
rect -3876 331076 -3276 331078
rect 587200 331076 587800 331078
rect -3876 330474 -3276 330476
rect 587200 330474 587800 330476
rect 0 327748 584000 330156
rect -1996 327428 -1396 327430
rect 585320 327428 585920 327430
rect -1996 326826 -1396 326828
rect 585320 326826 585920 326828
rect 0 320596 584000 326508
rect -8576 320276 -7976 320278
rect 591900 320276 592500 320278
rect -8576 319674 -7976 319676
rect 591900 319674 592500 319676
rect 0 316996 584000 319356
rect -6696 316676 -6096 316678
rect 590020 316676 590620 316678
rect -6696 316074 -6096 316076
rect 590020 316074 590620 316076
rect 0 313396 584000 315756
rect -4816 313076 -4216 313078
rect 588140 313076 588740 313078
rect -4816 312474 -4216 312476
rect 588140 312474 588740 312476
rect 0 309748 584000 312156
rect -2936 309428 -2336 309430
rect 586260 309428 586860 309430
rect -2936 308826 -2336 308828
rect 586260 308826 586860 308828
rect 0 302596 584000 308508
rect -7636 302276 -7036 302278
rect 590960 302276 591560 302278
rect -7636 301674 -7036 301676
rect 590960 301674 591560 301676
rect 0 298996 584000 301356
rect -5756 298676 -5156 298678
rect 589080 298676 589680 298678
rect -5756 298074 -5156 298076
rect 589080 298074 589680 298076
rect 0 295396 584000 297756
rect -3876 295076 -3276 295078
rect 587200 295076 587800 295078
rect -3876 294474 -3276 294476
rect 587200 294474 587800 294476
rect 0 291748 584000 294156
rect -1996 291428 -1396 291430
rect 585320 291428 585920 291430
rect -1996 290826 -1396 290828
rect 585320 290826 585920 290828
rect 0 284596 584000 290508
rect -8576 284276 -7976 284278
rect 591900 284276 592500 284278
rect -8576 283674 -7976 283676
rect 591900 283674 592500 283676
rect 0 280996 584000 283356
rect -6696 280676 -6096 280678
rect 590020 280676 590620 280678
rect -6696 280074 -6096 280076
rect 590020 280074 590620 280076
rect 0 277396 584000 279756
rect -4816 277076 -4216 277078
rect 588140 277076 588740 277078
rect -4816 276474 -4216 276476
rect 588140 276474 588740 276476
rect 0 273748 584000 276156
rect -2936 273428 -2336 273430
rect 586260 273428 586860 273430
rect -2936 272826 -2336 272828
rect 586260 272826 586860 272828
rect 0 266596 584000 272508
rect -7636 266276 -7036 266278
rect 590960 266276 591560 266278
rect -7636 265674 -7036 265676
rect 590960 265674 591560 265676
rect 0 262996 584000 265356
rect -5756 262676 -5156 262678
rect 589080 262676 589680 262678
rect -5756 262074 -5156 262076
rect 589080 262074 589680 262076
rect 0 259396 584000 261756
rect -3876 259076 -3276 259078
rect 587200 259076 587800 259078
rect -3876 258474 -3276 258476
rect 587200 258474 587800 258476
rect 0 255748 584000 258156
rect -1996 255428 -1396 255430
rect 585320 255428 585920 255430
rect -1996 254826 -1396 254828
rect 585320 254826 585920 254828
rect 0 248596 584000 254508
rect -8576 248276 -7976 248278
rect 591900 248276 592500 248278
rect -8576 247674 -7976 247676
rect 591900 247674 592500 247676
rect 0 244996 584000 247356
rect -6696 244676 -6096 244678
rect 590020 244676 590620 244678
rect -6696 244074 -6096 244076
rect 590020 244074 590620 244076
rect 0 241396 584000 243756
rect -4816 241076 -4216 241078
rect 588140 241076 588740 241078
rect -4816 240474 -4216 240476
rect 588140 240474 588740 240476
rect 0 237748 584000 240156
rect -2936 237428 -2336 237430
rect 586260 237428 586860 237430
rect -2936 236826 -2336 236828
rect 586260 236826 586860 236828
rect 0 230596 584000 236508
rect -7636 230276 -7036 230278
rect 590960 230276 591560 230278
rect -7636 229674 -7036 229676
rect 590960 229674 591560 229676
rect 0 226996 584000 229356
rect -5756 226676 -5156 226678
rect 589080 226676 589680 226678
rect -5756 226074 -5156 226076
rect 589080 226074 589680 226076
rect 0 223396 584000 225756
rect -3876 223076 -3276 223078
rect 587200 223076 587800 223078
rect -3876 222474 -3276 222476
rect 587200 222474 587800 222476
rect 0 219748 584000 222156
rect -1996 219428 -1396 219430
rect 585320 219428 585920 219430
rect -1996 218826 -1396 218828
rect 585320 218826 585920 218828
rect 0 212596 584000 218508
rect -8576 212276 -7976 212278
rect 591900 212276 592500 212278
rect -8576 211674 -7976 211676
rect 591900 211674 592500 211676
rect 0 208996 584000 211356
rect -6696 208676 -6096 208678
rect 590020 208676 590620 208678
rect -6696 208074 -6096 208076
rect 590020 208074 590620 208076
rect 0 205396 584000 207756
rect -4816 205076 -4216 205078
rect 588140 205076 588740 205078
rect -4816 204474 -4216 204476
rect 588140 204474 588740 204476
rect 0 201748 584000 204156
rect -2936 201428 -2336 201430
rect 586260 201428 586860 201430
rect -2936 200826 -2336 200828
rect 586260 200826 586860 200828
rect 0 194596 584000 200508
rect -7636 194276 -7036 194278
rect 590960 194276 591560 194278
rect -7636 193674 -7036 193676
rect 590960 193674 591560 193676
rect 0 190996 584000 193356
rect -5756 190676 -5156 190678
rect 589080 190676 589680 190678
rect -5756 190074 -5156 190076
rect 589080 190074 589680 190076
rect 0 187396 584000 189756
rect -3876 187076 -3276 187078
rect 587200 187076 587800 187078
rect -3876 186474 -3276 186476
rect 587200 186474 587800 186476
rect 0 183748 584000 186156
rect -1996 183428 -1396 183430
rect 585320 183428 585920 183430
rect -1996 182826 -1396 182828
rect 585320 182826 585920 182828
rect 0 176596 584000 182508
rect -8576 176276 -7976 176278
rect 591900 176276 592500 176278
rect -8576 175674 -7976 175676
rect 591900 175674 592500 175676
rect 0 172996 584000 175356
rect -6696 172676 -6096 172678
rect 590020 172676 590620 172678
rect -6696 172074 -6096 172076
rect 590020 172074 590620 172076
rect 0 169396 584000 171756
rect -4816 169076 -4216 169078
rect 588140 169076 588740 169078
rect -4816 168474 -4216 168476
rect 588140 168474 588740 168476
rect 0 165748 584000 168156
rect -2936 165428 -2336 165430
rect 586260 165428 586860 165430
rect -2936 164826 -2336 164828
rect 586260 164826 586860 164828
rect 0 158596 584000 164508
rect -7636 158276 -7036 158278
rect 590960 158276 591560 158278
rect -7636 157674 -7036 157676
rect 590960 157674 591560 157676
rect 0 154996 584000 157356
rect -5756 154676 -5156 154678
rect 589080 154676 589680 154678
rect -5756 154074 -5156 154076
rect 589080 154074 589680 154076
rect 0 151396 584000 153756
rect -3876 151076 -3276 151078
rect 587200 151076 587800 151078
rect -3876 150474 -3276 150476
rect 587200 150474 587800 150476
rect 0 147748 584000 150156
rect -1996 147428 -1396 147430
rect 585320 147428 585920 147430
rect -1996 146826 -1396 146828
rect 585320 146826 585920 146828
rect 0 140596 584000 146508
rect -8576 140276 -7976 140278
rect 591900 140276 592500 140278
rect -8576 139674 -7976 139676
rect 591900 139674 592500 139676
rect 0 136996 584000 139356
rect -6696 136676 -6096 136678
rect 590020 136676 590620 136678
rect -6696 136074 -6096 136076
rect 590020 136074 590620 136076
rect 0 133396 584000 135756
rect -4816 133076 -4216 133078
rect 588140 133076 588740 133078
rect -4816 132474 -4216 132476
rect 588140 132474 588740 132476
rect 0 129748 584000 132156
rect -2936 129428 -2336 129430
rect 586260 129428 586860 129430
rect -2936 128826 -2336 128828
rect 586260 128826 586860 128828
rect 0 122596 584000 128508
rect -7636 122276 -7036 122278
rect 590960 122276 591560 122278
rect -7636 121674 -7036 121676
rect 590960 121674 591560 121676
rect 0 118996 584000 121356
rect -5756 118676 -5156 118678
rect 589080 118676 589680 118678
rect -5756 118074 -5156 118076
rect 589080 118074 589680 118076
rect 0 115396 584000 117756
rect -3876 115076 -3276 115078
rect 587200 115076 587800 115078
rect -3876 114474 -3276 114476
rect 587200 114474 587800 114476
rect 0 111748 584000 114156
rect -1996 111428 -1396 111430
rect 585320 111428 585920 111430
rect -1996 110826 -1396 110828
rect 585320 110826 585920 110828
rect 0 104596 584000 110508
rect -8576 104276 -7976 104278
rect 591900 104276 592500 104278
rect -8576 103674 -7976 103676
rect 591900 103674 592500 103676
rect 0 100996 584000 103356
rect -6696 100676 -6096 100678
rect 590020 100676 590620 100678
rect -6696 100074 -6096 100076
rect 590020 100074 590620 100076
rect 0 97396 584000 99756
rect -4816 97076 -4216 97078
rect 588140 97076 588740 97078
rect -4816 96474 -4216 96476
rect 588140 96474 588740 96476
rect 0 93748 584000 96156
rect -2936 93428 -2336 93430
rect 586260 93428 586860 93430
rect -2936 92826 -2336 92828
rect 586260 92826 586860 92828
rect 0 86596 584000 92508
rect -7636 86276 -7036 86278
rect 590960 86276 591560 86278
rect -7636 85674 -7036 85676
rect 590960 85674 591560 85676
rect 0 82996 584000 85356
rect -5756 82676 -5156 82678
rect 589080 82676 589680 82678
rect -5756 82074 -5156 82076
rect 589080 82074 589680 82076
rect 0 79396 584000 81756
rect -3876 79076 -3276 79078
rect 587200 79076 587800 79078
rect -3876 78474 -3276 78476
rect 587200 78474 587800 78476
rect 0 75748 584000 78156
rect -1996 75428 -1396 75430
rect 585320 75428 585920 75430
rect -1996 74826 -1396 74828
rect 585320 74826 585920 74828
rect 0 68596 584000 74508
rect -8576 68276 -7976 68278
rect 591900 68276 592500 68278
rect -8576 67674 -7976 67676
rect 591900 67674 592500 67676
rect 0 64996 584000 67356
rect -6696 64676 -6096 64678
rect 590020 64676 590620 64678
rect -6696 64074 -6096 64076
rect 590020 64074 590620 64076
rect 0 61396 584000 63756
rect -4816 61076 -4216 61078
rect 588140 61076 588740 61078
rect -4816 60474 -4216 60476
rect 588140 60474 588740 60476
rect 0 57748 584000 60156
rect -2936 57428 -2336 57430
rect 586260 57428 586860 57430
rect -2936 56826 -2336 56828
rect 586260 56826 586860 56828
rect 0 50596 584000 56508
rect -7636 50276 -7036 50278
rect 590960 50276 591560 50278
rect -7636 49674 -7036 49676
rect 590960 49674 591560 49676
rect 0 46996 584000 49356
rect -5756 46676 -5156 46678
rect 589080 46676 589680 46678
rect -5756 46074 -5156 46076
rect 589080 46074 589680 46076
rect 0 43396 584000 45756
rect -3876 43076 -3276 43078
rect 587200 43076 587800 43078
rect -3876 42474 -3276 42476
rect 587200 42474 587800 42476
rect 0 39748 584000 42156
rect -1996 39428 -1396 39430
rect 585320 39428 585920 39430
rect -1996 38826 -1396 38828
rect 585320 38826 585920 38828
rect 0 32596 584000 38508
rect -8576 32276 -7976 32278
rect 591900 32276 592500 32278
rect -8576 31674 -7976 31676
rect 591900 31674 592500 31676
rect 0 28996 584000 31356
rect -6696 28676 -6096 28678
rect 590020 28676 590620 28678
rect -6696 28074 -6096 28076
rect 590020 28074 590620 28076
rect 0 25396 584000 27756
rect -4816 25076 -4216 25078
rect 588140 25076 588740 25078
rect -4816 24474 -4216 24476
rect 588140 24474 588740 24476
rect 0 21748 584000 24156
rect -2936 21428 -2336 21430
rect 586260 21428 586860 21430
rect -2936 20826 -2336 20828
rect 586260 20826 586860 20828
rect 0 14596 584000 20508
rect -7636 14276 -7036 14278
rect 590960 14276 591560 14278
rect -7636 13674 -7036 13676
rect 590960 13674 591560 13676
rect 0 10996 584000 13356
rect -5756 10676 -5156 10678
rect 589080 10676 589680 10678
rect -5756 10074 -5156 10076
rect 589080 10074 589680 10076
rect 0 7396 584000 9756
rect -3876 7076 -3276 7078
rect 587200 7076 587800 7078
rect -3876 6474 -3276 6476
rect 587200 6474 587800 6476
rect 0 3748 584000 6156
rect -1996 3428 -1396 3430
rect 585320 3428 585920 3430
rect -1996 2826 -1396 2828
rect 585320 2826 585920 2828
rect 0 0 584000 2508
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 532 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 541804 311388 542404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 505804 311388 506404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 469804 565820 470404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 433804 565820 434404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 397804 565820 398404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 253804 666052 254404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 217804 666052 218404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 181804 666052 182404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 145804 666052 146404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 109804 666052 110404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 73804 666052 74404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 37804 666052 38404 705800 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 469804 425812 470404 518048 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 433804 425812 434404 518048 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 397804 425812 398404 518048 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 518048 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 518048 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 518048 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 145804 495716 146404 518048 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 109804 495716 110404 518048 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 73804 495716 74404 518048 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 37804 495716 38404 518048 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 469804 311388 470404 358048 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 433804 311388 434404 358048 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 397804 311388 398404 358048 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 145804 325260 146404 358048 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 109804 325260 110404 358048 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 73804 325260 74404 358048 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 37804 325260 38404 358048 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 541804 208940 542404 238048 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 505804 208940 506404 238048 6 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 469804 208940 470404 238048 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 433804 208940 434404 238048 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 397804 208940 398404 238048 6 vccd1
port 678 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 238048 6 vccd1
port 679 nsew power bidirectional
rlabel metal4 s 109804 221452 110404 238048 6 vccd1
port 680 nsew power bidirectional
rlabel metal4 s 73804 221452 74404 238048 6 vccd1
port 681 nsew power bidirectional
rlabel metal4 s 37804 221452 38404 238048 6 vccd1
port 682 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 138048 6 vccd1
port 683 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 138048 6 vccd1
port 684 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 138048 6 vccd1
port 685 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 138048 6 vccd1
port 686 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 138048 6 vccd1
port 687 nsew power bidirectional
rlabel metal4 s 109804 111244 110404 138048 6 vccd1
port 688 nsew power bidirectional
rlabel metal4 s 73804 111244 74404 138048 6 vccd1
port 689 nsew power bidirectional
rlabel metal4 s 37804 111244 38404 138048 6 vccd1
port 690 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 18048 6 vccd1
port 691 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 18048 6 vccd1
port 692 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 18048 6 vccd1
port 693 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 694 nsew power bidirectional
rlabel metal5 s -2936 686828 586860 687428 6 vccd1
port 695 nsew power bidirectional
rlabel metal5 s -2936 650828 586860 651428 6 vccd1
port 696 nsew power bidirectional
rlabel metal5 s -2936 614828 586860 615428 6 vccd1
port 697 nsew power bidirectional
rlabel metal5 s -2936 578828 586860 579428 6 vccd1
port 698 nsew power bidirectional
rlabel metal5 s -2936 542828 586860 543428 6 vccd1
port 699 nsew power bidirectional
rlabel metal5 s -2936 506828 586860 507428 6 vccd1
port 700 nsew power bidirectional
rlabel metal5 s -2936 470828 586860 471428 6 vccd1
port 701 nsew power bidirectional
rlabel metal5 s -2936 434828 586860 435428 6 vccd1
port 702 nsew power bidirectional
rlabel metal5 s -2936 398828 586860 399428 6 vccd1
port 703 nsew power bidirectional
rlabel metal5 s -2936 362828 586860 363428 6 vccd1
port 704 nsew power bidirectional
rlabel metal5 s -2936 326828 586860 327428 6 vccd1
port 705 nsew power bidirectional
rlabel metal5 s -2936 290828 586860 291428 6 vccd1
port 706 nsew power bidirectional
rlabel metal5 s -2936 254828 586860 255428 6 vccd1
port 707 nsew power bidirectional
rlabel metal5 s -2936 218828 586860 219428 6 vccd1
port 708 nsew power bidirectional
rlabel metal5 s -2936 182828 586860 183428 6 vccd1
port 709 nsew power bidirectional
rlabel metal5 s -2936 146828 586860 147428 6 vccd1
port 710 nsew power bidirectional
rlabel metal5 s -2936 110828 586860 111428 6 vccd1
port 711 nsew power bidirectional
rlabel metal5 s -2936 74828 586860 75428 6 vccd1
port 712 nsew power bidirectional
rlabel metal5 s -2936 38828 586860 39428 6 vccd1
port 713 nsew power bidirectional
rlabel metal5 s -2936 2828 586860 3428 6 vccd1
port 714 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 715 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 559804 311388 560404 705800 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 523804 311388 524404 705800 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 487804 565820 488404 705800 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 451804 565820 452404 705800 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 415804 565820 416404 705800 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 705800 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 705800 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 705800 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 705800 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 235804 666052 236404 705800 6 vssd1
port 726 nsew ground bidirectional
rlabel metal4 s 199804 666052 200404 705800 6 vssd1
port 727 nsew ground bidirectional
rlabel metal4 s 163804 666052 164404 705800 6 vssd1
port 728 nsew ground bidirectional
rlabel metal4 s 127804 666052 128404 705800 6 vssd1
port 729 nsew ground bidirectional
rlabel metal4 s 91804 666052 92404 705800 6 vssd1
port 730 nsew ground bidirectional
rlabel metal4 s 55804 666052 56404 705800 6 vssd1
port 731 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 705800 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 733 nsew ground bidirectional
rlabel metal4 s 487804 425812 488404 518048 6 vssd1
port 734 nsew ground bidirectional
rlabel metal4 s 451804 425812 452404 518048 6 vssd1
port 735 nsew ground bidirectional
rlabel metal4 s 415804 425812 416404 518048 6 vssd1
port 736 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 518048 6 vssd1
port 737 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 518048 6 vssd1
port 738 nsew ground bidirectional
rlabel metal4 s 163804 495716 164404 518048 6 vssd1
port 739 nsew ground bidirectional
rlabel metal4 s 127804 495716 128404 518048 6 vssd1
port 740 nsew ground bidirectional
rlabel metal4 s 91804 495716 92404 518048 6 vssd1
port 741 nsew ground bidirectional
rlabel metal4 s 55804 495716 56404 518048 6 vssd1
port 742 nsew ground bidirectional
rlabel metal4 s 487804 311388 488404 358048 6 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 451804 311388 452404 358048 6 vssd1
port 744 nsew ground bidirectional
rlabel metal4 s 415804 311388 416404 358048 6 vssd1
port 745 nsew ground bidirectional
rlabel metal4 s 163804 325260 164404 358048 6 vssd1
port 746 nsew ground bidirectional
rlabel metal4 s 127804 325260 128404 358048 6 vssd1
port 747 nsew ground bidirectional
rlabel metal4 s 91804 325260 92404 358048 6 vssd1
port 748 nsew ground bidirectional
rlabel metal4 s 55804 325260 56404 358048 6 vssd1
port 749 nsew ground bidirectional
rlabel metal4 s 559804 208940 560404 238048 6 vssd1
port 750 nsew ground bidirectional
rlabel metal4 s 523804 208940 524404 238048 6 vssd1
port 751 nsew ground bidirectional
rlabel metal4 s 487804 208940 488404 238048 6 vssd1
port 752 nsew ground bidirectional
rlabel metal4 s 451804 208940 452404 238048 6 vssd1
port 753 nsew ground bidirectional
rlabel metal4 s 415804 208940 416404 238048 6 vssd1
port 754 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 238048 6 vssd1
port 755 nsew ground bidirectional
rlabel metal4 s 127804 221452 128404 238048 6 vssd1
port 756 nsew ground bidirectional
rlabel metal4 s 91804 221452 92404 238048 6 vssd1
port 757 nsew ground bidirectional
rlabel metal4 s 55804 221452 56404 238048 6 vssd1
port 758 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 138048 6 vssd1
port 759 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 138048 6 vssd1
port 760 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 138048 6 vssd1
port 761 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 138048 6 vssd1
port 762 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 138048 6 vssd1
port 763 nsew ground bidirectional
rlabel metal4 s 127804 111244 128404 138048 6 vssd1
port 764 nsew ground bidirectional
rlabel metal4 s 91804 111244 92404 138048 6 vssd1
port 765 nsew ground bidirectional
rlabel metal4 s 55804 111244 56404 138048 6 vssd1
port 766 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 18048 6 vssd1
port 767 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 18048 6 vssd1
port 768 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 18048 6 vssd1
port 769 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 770 nsew ground bidirectional
rlabel metal5 s -2936 668828 586860 669428 6 vssd1
port 771 nsew ground bidirectional
rlabel metal5 s -2936 632828 586860 633428 6 vssd1
port 772 nsew ground bidirectional
rlabel metal5 s -2936 596828 586860 597428 6 vssd1
port 773 nsew ground bidirectional
rlabel metal5 s -2936 560828 586860 561428 6 vssd1
port 774 nsew ground bidirectional
rlabel metal5 s -2936 524828 586860 525428 6 vssd1
port 775 nsew ground bidirectional
rlabel metal5 s -2936 488828 586860 489428 6 vssd1
port 776 nsew ground bidirectional
rlabel metal5 s -2936 452828 586860 453428 6 vssd1
port 777 nsew ground bidirectional
rlabel metal5 s -2936 416828 586860 417428 6 vssd1
port 778 nsew ground bidirectional
rlabel metal5 s -2936 380828 586860 381428 6 vssd1
port 779 nsew ground bidirectional
rlabel metal5 s -2936 344828 586860 345428 6 vssd1
port 780 nsew ground bidirectional
rlabel metal5 s -2936 308828 586860 309428 6 vssd1
port 781 nsew ground bidirectional
rlabel metal5 s -2936 272828 586860 273428 6 vssd1
port 782 nsew ground bidirectional
rlabel metal5 s -2936 236828 586860 237428 6 vssd1
port 783 nsew ground bidirectional
rlabel metal5 s -2936 200828 586860 201428 6 vssd1
port 784 nsew ground bidirectional
rlabel metal5 s -2936 164828 586860 165428 6 vssd1
port 785 nsew ground bidirectional
rlabel metal5 s -2936 128828 586860 129428 6 vssd1
port 786 nsew ground bidirectional
rlabel metal5 s -2936 92828 586860 93428 6 vssd1
port 787 nsew ground bidirectional
rlabel metal5 s -2936 56828 586860 57428 6 vssd1
port 788 nsew ground bidirectional
rlabel metal5 s -2936 20828 586860 21428 6 vssd1
port 789 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 790 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 791 nsew power bidirectional
rlabel metal4 s 545404 311436 546004 707680 6 vccd2
port 792 nsew power bidirectional
rlabel metal4 s 509404 311436 510004 707680 6 vccd2
port 793 nsew power bidirectional
rlabel metal4 s 473404 565868 474004 707680 6 vccd2
port 794 nsew power bidirectional
rlabel metal4 s 437404 565868 438004 707680 6 vccd2
port 795 nsew power bidirectional
rlabel metal4 s 401404 565868 402004 707680 6 vccd2
port 796 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 707680 6 vccd2
port 797 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 707680 6 vccd2
port 798 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 707680 6 vccd2
port 799 nsew power bidirectional
rlabel metal4 s 257404 666100 258004 707680 6 vccd2
port 800 nsew power bidirectional
rlabel metal4 s 221404 666100 222004 707680 6 vccd2
port 801 nsew power bidirectional
rlabel metal4 s 185404 666100 186004 707680 6 vccd2
port 802 nsew power bidirectional
rlabel metal4 s 149404 666100 150004 707680 6 vccd2
port 803 nsew power bidirectional
rlabel metal4 s 113404 666100 114004 707680 6 vccd2
port 804 nsew power bidirectional
rlabel metal4 s 77404 666100 78004 707680 6 vccd2
port 805 nsew power bidirectional
rlabel metal4 s 41404 666100 42004 707680 6 vccd2
port 806 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 807 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 808 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 809 nsew power bidirectional
rlabel metal4 s 473404 425860 474004 518000 6 vccd2
port 810 nsew power bidirectional
rlabel metal4 s 437404 425860 438004 518000 6 vccd2
port 811 nsew power bidirectional
rlabel metal4 s 401404 425860 402004 518000 6 vccd2
port 812 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 518000 6 vccd2
port 813 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 518000 6 vccd2
port 814 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 518000 6 vccd2
port 815 nsew power bidirectional
rlabel metal4 s 149404 495764 150004 518000 6 vccd2
port 816 nsew power bidirectional
rlabel metal4 s 113404 495764 114004 518000 6 vccd2
port 817 nsew power bidirectional
rlabel metal4 s 77404 495764 78004 518000 6 vccd2
port 818 nsew power bidirectional
rlabel metal4 s 41404 495764 42004 518000 6 vccd2
port 819 nsew power bidirectional
rlabel metal4 s 473404 311436 474004 358000 6 vccd2
port 820 nsew power bidirectional
rlabel metal4 s 437404 311436 438004 358000 6 vccd2
port 821 nsew power bidirectional
rlabel metal4 s 401404 311436 402004 358000 6 vccd2
port 822 nsew power bidirectional
rlabel metal4 s 149404 325308 150004 358000 6 vccd2
port 823 nsew power bidirectional
rlabel metal4 s 113404 325308 114004 358000 6 vccd2
port 824 nsew power bidirectional
rlabel metal4 s 77404 325308 78004 358000 6 vccd2
port 825 nsew power bidirectional
rlabel metal4 s 41404 325308 42004 358000 6 vccd2
port 826 nsew power bidirectional
rlabel metal4 s 545404 208988 546004 238000 6 vccd2
port 827 nsew power bidirectional
rlabel metal4 s 509404 208988 510004 238000 6 vccd2
port 828 nsew power bidirectional
rlabel metal4 s 473404 208988 474004 238000 6 vccd2
port 829 nsew power bidirectional
rlabel metal4 s 437404 208988 438004 238000 6 vccd2
port 830 nsew power bidirectional
rlabel metal4 s 401404 208988 402004 238000 6 vccd2
port 831 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 238000 6 vccd2
port 832 nsew power bidirectional
rlabel metal4 s 113404 221500 114004 238000 6 vccd2
port 833 nsew power bidirectional
rlabel metal4 s 77404 221500 78004 238000 6 vccd2
port 834 nsew power bidirectional
rlabel metal4 s 41404 221500 42004 238000 6 vccd2
port 835 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 138000 6 vccd2
port 836 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 138000 6 vccd2
port 837 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 138000 6 vccd2
port 838 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 138000 6 vccd2
port 839 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 138000 6 vccd2
port 840 nsew power bidirectional
rlabel metal4 s 113404 111292 114004 138000 6 vccd2
port 841 nsew power bidirectional
rlabel metal4 s 77404 111292 78004 138000 6 vccd2
port 842 nsew power bidirectional
rlabel metal4 s 41404 111292 42004 138000 6 vccd2
port 843 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 18000 6 vccd2
port 844 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 18000 6 vccd2
port 845 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 18000 6 vccd2
port 846 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 847 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 848 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 849 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 850 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 851 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 852 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 853 nsew power bidirectional
rlabel metal5 s -4816 474476 588740 475076 6 vccd2
port 854 nsew power bidirectional
rlabel metal5 s -4816 438476 588740 439076 6 vccd2
port 855 nsew power bidirectional
rlabel metal5 s -4816 402476 588740 403076 6 vccd2
port 856 nsew power bidirectional
rlabel metal5 s -4816 366476 588740 367076 6 vccd2
port 857 nsew power bidirectional
rlabel metal5 s -4816 330476 588740 331076 6 vccd2
port 858 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 859 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 860 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 861 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 862 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 863 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 864 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 865 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 866 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 867 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 868 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 869 nsew ground bidirectional
rlabel metal4 s 563404 208988 564004 707680 6 vssd2
port 870 nsew ground bidirectional
rlabel metal4 s 527404 311436 528004 707680 6 vssd2
port 871 nsew ground bidirectional
rlabel metal4 s 491404 565868 492004 707680 6 vssd2
port 872 nsew ground bidirectional
rlabel metal4 s 455404 565868 456004 707680 6 vssd2
port 873 nsew ground bidirectional
rlabel metal4 s 419404 565868 420004 707680 6 vssd2
port 874 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 707680 6 vssd2
port 875 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 707680 6 vssd2
port 876 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 707680 6 vssd2
port 877 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 707680 6 vssd2
port 878 nsew ground bidirectional
rlabel metal4 s 239404 666100 240004 707680 6 vssd2
port 879 nsew ground bidirectional
rlabel metal4 s 203404 666100 204004 707680 6 vssd2
port 880 nsew ground bidirectional
rlabel metal4 s 167404 666100 168004 707680 6 vssd2
port 881 nsew ground bidirectional
rlabel metal4 s 131404 666100 132004 707680 6 vssd2
port 882 nsew ground bidirectional
rlabel metal4 s 95404 666100 96004 707680 6 vssd2
port 883 nsew ground bidirectional
rlabel metal4 s 59404 666100 60004 707680 6 vssd2
port 884 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2
port 885 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 886 nsew ground bidirectional
rlabel metal4 s 491404 425860 492004 518000 6 vssd2
port 887 nsew ground bidirectional
rlabel metal4 s 455404 425860 456004 518000 6 vssd2
port 888 nsew ground bidirectional
rlabel metal4 s 419404 425860 420004 518000 6 vssd2
port 889 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 518000 6 vssd2
port 890 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 518000 6 vssd2
port 891 nsew ground bidirectional
rlabel metal4 s 167404 495764 168004 518000 6 vssd2
port 892 nsew ground bidirectional
rlabel metal4 s 131404 495764 132004 518000 6 vssd2
port 893 nsew ground bidirectional
rlabel metal4 s 95404 495764 96004 518000 6 vssd2
port 894 nsew ground bidirectional
rlabel metal4 s 59404 495764 60004 518000 6 vssd2
port 895 nsew ground bidirectional
rlabel metal4 s 491404 311436 492004 358000 6 vssd2
port 896 nsew ground bidirectional
rlabel metal4 s 455404 311436 456004 358000 6 vssd2
port 897 nsew ground bidirectional
rlabel metal4 s 419404 311436 420004 358000 6 vssd2
port 898 nsew ground bidirectional
rlabel metal4 s 167404 325308 168004 358000 6 vssd2
port 899 nsew ground bidirectional
rlabel metal4 s 131404 325308 132004 358000 6 vssd2
port 900 nsew ground bidirectional
rlabel metal4 s 95404 325308 96004 358000 6 vssd2
port 901 nsew ground bidirectional
rlabel metal4 s 59404 325308 60004 358000 6 vssd2
port 902 nsew ground bidirectional
rlabel metal4 s 527404 208988 528004 238000 6 vssd2
port 903 nsew ground bidirectional
rlabel metal4 s 491404 208988 492004 238000 6 vssd2
port 904 nsew ground bidirectional
rlabel metal4 s 455404 208988 456004 238000 6 vssd2
port 905 nsew ground bidirectional
rlabel metal4 s 419404 208988 420004 238000 6 vssd2
port 906 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 238000 6 vssd2
port 907 nsew ground bidirectional
rlabel metal4 s 131404 221500 132004 238000 6 vssd2
port 908 nsew ground bidirectional
rlabel metal4 s 95404 221500 96004 238000 6 vssd2
port 909 nsew ground bidirectional
rlabel metal4 s 59404 221500 60004 238000 6 vssd2
port 910 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 138000 6 vssd2
port 911 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 138000 6 vssd2
port 912 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 138000 6 vssd2
port 913 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 138000 6 vssd2
port 914 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 138000 6 vssd2
port 915 nsew ground bidirectional
rlabel metal4 s 131404 111292 132004 138000 6 vssd2
port 916 nsew ground bidirectional
rlabel metal4 s 95404 111292 96004 138000 6 vssd2
port 917 nsew ground bidirectional
rlabel metal4 s 59404 111292 60004 138000 6 vssd2
port 918 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 18000 6 vssd2
port 919 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 18000 6 vssd2
port 920 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 18000 6 vssd2
port 921 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 922 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 923 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 924 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 925 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 926 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 927 nsew ground bidirectional
rlabel metal5 s -4816 492476 588740 493076 6 vssd2
port 928 nsew ground bidirectional
rlabel metal5 s -4816 456476 588740 457076 6 vssd2
port 929 nsew ground bidirectional
rlabel metal5 s -4816 420476 588740 421076 6 vssd2
port 930 nsew ground bidirectional
rlabel metal5 s -4816 384476 588740 385076 6 vssd2
port 931 nsew ground bidirectional
rlabel metal5 s -4816 348476 588740 349076 6 vssd2
port 932 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 933 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 934 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 935 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 936 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 937 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 938 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 939 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 940 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 941 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 942 nsew ground bidirectional
rlabel metal4 s 549004 311436 549604 709560 6 vdda1
port 943 nsew power bidirectional
rlabel metal4 s 513004 311436 513604 709560 6 vdda1
port 944 nsew power bidirectional
rlabel metal4 s 477004 565868 477604 709560 6 vdda1
port 945 nsew power bidirectional
rlabel metal4 s 441004 565868 441604 709560 6 vdda1
port 946 nsew power bidirectional
rlabel metal4 s 405004 565868 405604 709560 6 vdda1
port 947 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 709560 6 vdda1
port 948 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 709560 6 vdda1
port 949 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 709560 6 vdda1
port 950 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 709560 6 vdda1
port 951 nsew power bidirectional
rlabel metal4 s 225004 666100 225604 709560 6 vdda1
port 952 nsew power bidirectional
rlabel metal4 s 189004 666100 189604 709560 6 vdda1
port 953 nsew power bidirectional
rlabel metal4 s 153004 666100 153604 709560 6 vdda1
port 954 nsew power bidirectional
rlabel metal4 s 117004 666100 117604 709560 6 vdda1
port 955 nsew power bidirectional
rlabel metal4 s 81004 666100 81604 709560 6 vdda1
port 956 nsew power bidirectional
rlabel metal4 s 45004 666100 45604 709560 6 vdda1
port 957 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 958 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 959 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 960 nsew power bidirectional
rlabel metal4 s 477004 425860 477604 518000 6 vdda1
port 961 nsew power bidirectional
rlabel metal4 s 441004 425860 441604 518000 6 vdda1
port 962 nsew power bidirectional
rlabel metal4 s 405004 425860 405604 518000 6 vdda1
port 963 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 518000 6 vdda1
port 964 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 518000 6 vdda1
port 965 nsew power bidirectional
rlabel metal4 s 153004 495764 153604 518000 6 vdda1
port 966 nsew power bidirectional
rlabel metal4 s 117004 495764 117604 518000 6 vdda1
port 967 nsew power bidirectional
rlabel metal4 s 81004 495764 81604 518000 6 vdda1
port 968 nsew power bidirectional
rlabel metal4 s 45004 495764 45604 518000 6 vdda1
port 969 nsew power bidirectional
rlabel metal4 s 477004 311436 477604 358000 6 vdda1
port 970 nsew power bidirectional
rlabel metal4 s 441004 311436 441604 358000 6 vdda1
port 971 nsew power bidirectional
rlabel metal4 s 405004 311436 405604 358000 6 vdda1
port 972 nsew power bidirectional
rlabel metal4 s 153004 325308 153604 358000 6 vdda1
port 973 nsew power bidirectional
rlabel metal4 s 117004 325308 117604 358000 6 vdda1
port 974 nsew power bidirectional
rlabel metal4 s 81004 325308 81604 358000 6 vdda1
port 975 nsew power bidirectional
rlabel metal4 s 45004 325308 45604 358000 6 vdda1
port 976 nsew power bidirectional
rlabel metal4 s 549004 208988 549604 238000 6 vdda1
port 977 nsew power bidirectional
rlabel metal4 s 513004 208988 513604 238000 6 vdda1
port 978 nsew power bidirectional
rlabel metal4 s 477004 208988 477604 238000 6 vdda1
port 979 nsew power bidirectional
rlabel metal4 s 441004 208988 441604 238000 6 vdda1
port 980 nsew power bidirectional
rlabel metal4 s 405004 208988 405604 238000 6 vdda1
port 981 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 238000 6 vdda1
port 982 nsew power bidirectional
rlabel metal4 s 117004 221500 117604 238000 6 vdda1
port 983 nsew power bidirectional
rlabel metal4 s 81004 221500 81604 238000 6 vdda1
port 984 nsew power bidirectional
rlabel metal4 s 45004 221500 45604 238000 6 vdda1
port 985 nsew power bidirectional
rlabel metal4 s 549004 -5624 549604 138000 6 vdda1
port 986 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 138000 6 vdda1
port 987 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 138000 6 vdda1
port 988 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 138000 6 vdda1
port 989 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 138000 6 vdda1
port 990 nsew power bidirectional
rlabel metal4 s 117004 111292 117604 138000 6 vdda1
port 991 nsew power bidirectional
rlabel metal4 s 81004 111292 81604 138000 6 vdda1
port 992 nsew power bidirectional
rlabel metal4 s 45004 111292 45604 138000 6 vdda1
port 993 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 18000 6 vdda1
port 994 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 18000 6 vdda1
port 995 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 18000 6 vdda1
port 996 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 997 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 998 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 999 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 1000 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 1001 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 1002 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 1003 nsew power bidirectional
rlabel metal5 s -6696 478076 590620 478676 6 vdda1
port 1004 nsew power bidirectional
rlabel metal5 s -6696 442076 590620 442676 6 vdda1
port 1005 nsew power bidirectional
rlabel metal5 s -6696 406076 590620 406676 6 vdda1
port 1006 nsew power bidirectional
rlabel metal5 s -6696 370076 590620 370676 6 vdda1
port 1007 nsew power bidirectional
rlabel metal5 s -6696 334076 590620 334676 6 vdda1
port 1008 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 1009 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 1010 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 1011 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 1012 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 1013 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 1014 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 1015 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 1016 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 1017 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 1018 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 1019 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1
port 1020 nsew ground bidirectional
rlabel metal4 s 531004 311436 531604 709560 6 vssa1
port 1021 nsew ground bidirectional
rlabel metal4 s 495004 565868 495604 709560 6 vssa1
port 1022 nsew ground bidirectional
rlabel metal4 s 459004 565868 459604 709560 6 vssa1
port 1023 nsew ground bidirectional
rlabel metal4 s 423004 565868 423604 709560 6 vssa1
port 1024 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 709560 6 vssa1
port 1025 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 709560 6 vssa1
port 1026 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 709560 6 vssa1
port 1027 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 709560 6 vssa1
port 1028 nsew ground bidirectional
rlabel metal4 s 243004 666100 243604 709560 6 vssa1
port 1029 nsew ground bidirectional
rlabel metal4 s 207004 666100 207604 709560 6 vssa1
port 1030 nsew ground bidirectional
rlabel metal4 s 171004 666100 171604 709560 6 vssa1
port 1031 nsew ground bidirectional
rlabel metal4 s 135004 666100 135604 709560 6 vssa1
port 1032 nsew ground bidirectional
rlabel metal4 s 99004 666100 99604 709560 6 vssa1
port 1033 nsew ground bidirectional
rlabel metal4 s 63004 666100 63604 709560 6 vssa1
port 1034 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1
port 1035 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 1036 nsew ground bidirectional
rlabel metal4 s 495004 425860 495604 518000 6 vssa1
port 1037 nsew ground bidirectional
rlabel metal4 s 459004 425860 459604 518000 6 vssa1
port 1038 nsew ground bidirectional
rlabel metal4 s 423004 425860 423604 518000 6 vssa1
port 1039 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 518000 6 vssa1
port 1040 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 518000 6 vssa1
port 1041 nsew ground bidirectional
rlabel metal4 s 171004 495764 171604 518000 6 vssa1
port 1042 nsew ground bidirectional
rlabel metal4 s 135004 495764 135604 518000 6 vssa1
port 1043 nsew ground bidirectional
rlabel metal4 s 99004 495764 99604 518000 6 vssa1
port 1044 nsew ground bidirectional
rlabel metal4 s 63004 495764 63604 518000 6 vssa1
port 1045 nsew ground bidirectional
rlabel metal4 s 495004 311436 495604 358000 6 vssa1
port 1046 nsew ground bidirectional
rlabel metal4 s 459004 311436 459604 358000 6 vssa1
port 1047 nsew ground bidirectional
rlabel metal4 s 423004 311436 423604 358000 6 vssa1
port 1048 nsew ground bidirectional
rlabel metal4 s 171004 325308 171604 358000 6 vssa1
port 1049 nsew ground bidirectional
rlabel metal4 s 135004 325308 135604 358000 6 vssa1
port 1050 nsew ground bidirectional
rlabel metal4 s 99004 325308 99604 358000 6 vssa1
port 1051 nsew ground bidirectional
rlabel metal4 s 63004 325308 63604 358000 6 vssa1
port 1052 nsew ground bidirectional
rlabel metal4 s 531004 208988 531604 238000 6 vssa1
port 1053 nsew ground bidirectional
rlabel metal4 s 495004 208988 495604 238000 6 vssa1
port 1054 nsew ground bidirectional
rlabel metal4 s 459004 208988 459604 238000 6 vssa1
port 1055 nsew ground bidirectional
rlabel metal4 s 423004 208988 423604 238000 6 vssa1
port 1056 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 238000 6 vssa1
port 1057 nsew ground bidirectional
rlabel metal4 s 135004 221500 135604 238000 6 vssa1
port 1058 nsew ground bidirectional
rlabel metal4 s 99004 221500 99604 238000 6 vssa1
port 1059 nsew ground bidirectional
rlabel metal4 s 63004 221500 63604 238000 6 vssa1
port 1060 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 138000 6 vssa1
port 1061 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 138000 6 vssa1
port 1062 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 138000 6 vssa1
port 1063 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 138000 6 vssa1
port 1064 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 138000 6 vssa1
port 1065 nsew ground bidirectional
rlabel metal4 s 99004 111292 99604 138000 6 vssa1
port 1066 nsew ground bidirectional
rlabel metal4 s 63004 111292 63604 138000 6 vssa1
port 1067 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 18000 6 vssa1
port 1068 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 18000 6 vssa1
port 1069 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 1070 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 1071 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 1072 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 1073 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 1074 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 1075 nsew ground bidirectional
rlabel metal5 s -6696 496076 590620 496676 6 vssa1
port 1076 nsew ground bidirectional
rlabel metal5 s -6696 460076 590620 460676 6 vssa1
port 1077 nsew ground bidirectional
rlabel metal5 s -6696 424076 590620 424676 6 vssa1
port 1078 nsew ground bidirectional
rlabel metal5 s -6696 388076 590620 388676 6 vssa1
port 1079 nsew ground bidirectional
rlabel metal5 s -6696 352076 590620 352676 6 vssa1
port 1080 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 1081 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 1082 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 1083 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 1084 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 1085 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 1086 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 1087 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 1088 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 1089 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 1090 nsew ground bidirectional
rlabel metal4 s 552604 311436 553204 711440 6 vdda2
port 1091 nsew power bidirectional
rlabel metal4 s 516604 311436 517204 711440 6 vdda2
port 1092 nsew power bidirectional
rlabel metal4 s 480604 565868 481204 711440 6 vdda2
port 1093 nsew power bidirectional
rlabel metal4 s 444604 565868 445204 711440 6 vdda2
port 1094 nsew power bidirectional
rlabel metal4 s 408604 565868 409204 711440 6 vdda2
port 1095 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 711440 6 vdda2
port 1096 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 711440 6 vdda2
port 1097 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 711440 6 vdda2
port 1098 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 711440 6 vdda2
port 1099 nsew power bidirectional
rlabel metal4 s 228604 666100 229204 711440 6 vdda2
port 1100 nsew power bidirectional
rlabel metal4 s 192604 666100 193204 711440 6 vdda2
port 1101 nsew power bidirectional
rlabel metal4 s 156604 666100 157204 711440 6 vdda2
port 1102 nsew power bidirectional
rlabel metal4 s 120604 666100 121204 711440 6 vdda2
port 1103 nsew power bidirectional
rlabel metal4 s 84604 666100 85204 711440 6 vdda2
port 1104 nsew power bidirectional
rlabel metal4 s 48604 666100 49204 711440 6 vdda2
port 1105 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 1106 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 1107 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 1108 nsew power bidirectional
rlabel metal4 s 480604 425860 481204 518000 6 vdda2
port 1109 nsew power bidirectional
rlabel metal4 s 444604 425860 445204 518000 6 vdda2
port 1110 nsew power bidirectional
rlabel metal4 s 408604 425860 409204 518000 6 vdda2
port 1111 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 518000 6 vdda2
port 1112 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 518000 6 vdda2
port 1113 nsew power bidirectional
rlabel metal4 s 156604 495764 157204 518000 6 vdda2
port 1114 nsew power bidirectional
rlabel metal4 s 120604 495764 121204 518000 6 vdda2
port 1115 nsew power bidirectional
rlabel metal4 s 84604 495764 85204 518000 6 vdda2
port 1116 nsew power bidirectional
rlabel metal4 s 48604 495764 49204 518000 6 vdda2
port 1117 nsew power bidirectional
rlabel metal4 s 480604 311436 481204 358000 6 vdda2
port 1118 nsew power bidirectional
rlabel metal4 s 444604 311436 445204 358000 6 vdda2
port 1119 nsew power bidirectional
rlabel metal4 s 408604 311436 409204 358000 6 vdda2
port 1120 nsew power bidirectional
rlabel metal4 s 156604 325308 157204 358000 6 vdda2
port 1121 nsew power bidirectional
rlabel metal4 s 120604 325308 121204 358000 6 vdda2
port 1122 nsew power bidirectional
rlabel metal4 s 84604 325308 85204 358000 6 vdda2
port 1123 nsew power bidirectional
rlabel metal4 s 48604 325308 49204 358000 6 vdda2
port 1124 nsew power bidirectional
rlabel metal4 s 552604 208988 553204 238000 6 vdda2
port 1125 nsew power bidirectional
rlabel metal4 s 516604 208988 517204 238000 6 vdda2
port 1126 nsew power bidirectional
rlabel metal4 s 480604 208988 481204 238000 6 vdda2
port 1127 nsew power bidirectional
rlabel metal4 s 444604 208988 445204 238000 6 vdda2
port 1128 nsew power bidirectional
rlabel metal4 s 408604 208988 409204 238000 6 vdda2
port 1129 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 238000 6 vdda2
port 1130 nsew power bidirectional
rlabel metal4 s 120604 221500 121204 238000 6 vdda2
port 1131 nsew power bidirectional
rlabel metal4 s 84604 221500 85204 238000 6 vdda2
port 1132 nsew power bidirectional
rlabel metal4 s 48604 221500 49204 238000 6 vdda2
port 1133 nsew power bidirectional
rlabel metal4 s 552604 -7504 553204 138000 6 vdda2
port 1134 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 138000 6 vdda2
port 1135 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 138000 6 vdda2
port 1136 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 138000 6 vdda2
port 1137 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 138000 6 vdda2
port 1138 nsew power bidirectional
rlabel metal4 s 120604 111292 121204 138000 6 vdda2
port 1139 nsew power bidirectional
rlabel metal4 s 84604 111292 85204 138000 6 vdda2
port 1140 nsew power bidirectional
rlabel metal4 s 48604 111292 49204 138000 6 vdda2
port 1141 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 18000 6 vdda2
port 1142 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 18000 6 vdda2
port 1143 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 18000 6 vdda2
port 1144 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1145 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 1146 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 1147 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 1148 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 1149 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 1150 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 1151 nsew power bidirectional
rlabel metal5 s -8576 481676 592500 482276 6 vdda2
port 1152 nsew power bidirectional
rlabel metal5 s -8576 445676 592500 446276 6 vdda2
port 1153 nsew power bidirectional
rlabel metal5 s -8576 409676 592500 410276 6 vdda2
port 1154 nsew power bidirectional
rlabel metal5 s -8576 373676 592500 374276 6 vdda2
port 1155 nsew power bidirectional
rlabel metal5 s -8576 337676 592500 338276 6 vdda2
port 1156 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 1157 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 1158 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 1159 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 1160 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 1161 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 1162 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 1163 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 1164 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 1165 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1166 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1167 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2
port 1168 nsew ground bidirectional
rlabel metal4 s 534604 311436 535204 711440 6 vssa2
port 1169 nsew ground bidirectional
rlabel metal4 s 498604 311436 499204 711440 6 vssa2
port 1170 nsew ground bidirectional
rlabel metal4 s 462604 565868 463204 711440 6 vssa2
port 1171 nsew ground bidirectional
rlabel metal4 s 426604 565868 427204 711440 6 vssa2
port 1172 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 711440 6 vssa2
port 1173 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 711440 6 vssa2
port 1174 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 711440 6 vssa2
port 1175 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 711440 6 vssa2
port 1176 nsew ground bidirectional
rlabel metal4 s 246604 666100 247204 711440 6 vssa2
port 1177 nsew ground bidirectional
rlabel metal4 s 210604 666100 211204 711440 6 vssa2
port 1178 nsew ground bidirectional
rlabel metal4 s 174604 666100 175204 711440 6 vssa2
port 1179 nsew ground bidirectional
rlabel metal4 s 138604 666100 139204 711440 6 vssa2
port 1180 nsew ground bidirectional
rlabel metal4 s 102604 666100 103204 711440 6 vssa2
port 1181 nsew ground bidirectional
rlabel metal4 s 66604 666100 67204 711440 6 vssa2
port 1182 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2
port 1183 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1184 nsew ground bidirectional
rlabel metal4 s 462604 425860 463204 518000 6 vssa2
port 1185 nsew ground bidirectional
rlabel metal4 s 426604 425860 427204 518000 6 vssa2
port 1186 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 518000 6 vssa2
port 1187 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 518000 6 vssa2
port 1188 nsew ground bidirectional
rlabel metal4 s 174604 495764 175204 518000 6 vssa2
port 1189 nsew ground bidirectional
rlabel metal4 s 138604 495764 139204 518000 6 vssa2
port 1190 nsew ground bidirectional
rlabel metal4 s 102604 495764 103204 518000 6 vssa2
port 1191 nsew ground bidirectional
rlabel metal4 s 66604 495764 67204 518000 6 vssa2
port 1192 nsew ground bidirectional
rlabel metal4 s 462604 311436 463204 358000 6 vssa2
port 1193 nsew ground bidirectional
rlabel metal4 s 426604 311436 427204 358000 6 vssa2
port 1194 nsew ground bidirectional
rlabel metal4 s 174604 325308 175204 358000 6 vssa2
port 1195 nsew ground bidirectional
rlabel metal4 s 138604 325308 139204 358000 6 vssa2
port 1196 nsew ground bidirectional
rlabel metal4 s 102604 325308 103204 358000 6 vssa2
port 1197 nsew ground bidirectional
rlabel metal4 s 66604 325308 67204 358000 6 vssa2
port 1198 nsew ground bidirectional
rlabel metal4 s 534604 208988 535204 238000 6 vssa2
port 1199 nsew ground bidirectional
rlabel metal4 s 498604 208988 499204 238000 6 vssa2
port 1200 nsew ground bidirectional
rlabel metal4 s 462604 208988 463204 238000 6 vssa2
port 1201 nsew ground bidirectional
rlabel metal4 s 426604 208988 427204 238000 6 vssa2
port 1202 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 238000 6 vssa2
port 1203 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 238000 6 vssa2
port 1204 nsew ground bidirectional
rlabel metal4 s 102604 221500 103204 238000 6 vssa2
port 1205 nsew ground bidirectional
rlabel metal4 s 66604 221500 67204 238000 6 vssa2
port 1206 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 138000 6 vssa2
port 1207 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 138000 6 vssa2
port 1208 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 138000 6 vssa2
port 1209 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 138000 6 vssa2
port 1210 nsew ground bidirectional
rlabel metal4 s 102604 111292 103204 138000 6 vssa2
port 1211 nsew ground bidirectional
rlabel metal4 s 66604 111292 67204 138000 6 vssa2
port 1212 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 18000 6 vssa2
port 1213 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 18000 6 vssa2
port 1214 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1215 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 1216 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 1217 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 1218 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 1219 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 1220 nsew ground bidirectional
rlabel metal5 s -8576 499676 592500 500276 6 vssa2
port 1221 nsew ground bidirectional
rlabel metal5 s -8576 463676 592500 464276 6 vssa2
port 1222 nsew ground bidirectional
rlabel metal5 s -8576 427676 592500 428276 6 vssa2
port 1223 nsew ground bidirectional
rlabel metal5 s -8576 391676 592500 392276 6 vssa2
port 1224 nsew ground bidirectional
rlabel metal5 s -8576 355676 592500 356276 6 vssa2
port 1225 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 1226 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 1227 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 1228 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 1229 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 1230 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 1231 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 1232 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 1233 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 1234 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1235 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 123075158
string GDS_START 36877760
<< end >>

