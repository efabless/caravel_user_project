`default_nettype none
//-----------------------------------------------------
// Project Name : Register File
// Function     : Rergiter bank data 
// Description  : This is the main processor
// Coder        : Ivan Rodriguez Ferrandez  AND Alvaro Jover-Alvarez

//***Headers***

//***Module***
module register_data #(
        parameter integer WORD_SIZE = 32,
        parameter integer REGISTERS = 32,
        parameter integer REGDIRSIZE = 5,
        parameter integer ECCBITS = 7,
        parameter integer WHISBONE_ADR = 32,
        parameter [31:0]  ADDRBASE     = 32'h3000_0000,
        parameter [31:0]  REGISTERDATA  = ADDRBASE
    )
    (
        input  clk_i,
        input  rst_i ,
        input  [WORD_SIZE + ECCBITS - 1 : 0] data_to_register_i ,
        input  [REGDIRSIZE - 1 : 0] register_i ,
        input  [WHISBONE_ADR - 1 : 0] whisbone_addr_i,
        input  wregister_i ,
        input  rregister_i ,
        input  valid_i, 
        input  [3 : 0] wstrb_i,
        input  [WORD_SIZE -1 : 0] wdata_i,
        input  wbs_we_i,
        output reg [WORD_SIZE + ECCBITS -1: 0] store_data_o ,
        output reg ready_o,
        output reg [WORD_SIZE - 1 : 0] rdata_o
    );

//***Internal logic generated by compiler***  


//***Dumped Internal logic***
    // register bank
    reg [WORD_SIZE + ECCBITS -1:0] r[0:REGISTERS-1];
    wire [ECCBITS - 1:0] parity_bits;

    //request

    always @(*) begin
        // calculate last parity bit
        if (rst_i) begin

            r[0] = {WORD_SIZE + ECCBITS{1'b0}};
            r[1] = {WORD_SIZE + ECCBITS{1'b0}};
            r[2] = {WORD_SIZE + ECCBITS{1'b0}};
            r[3] = {WORD_SIZE + ECCBITS{1'b0}};
            r[4] = {WORD_SIZE + ECCBITS{1'b0}};
            r[5] = {WORD_SIZE + ECCBITS{1'b0}};
            r[6] = {WORD_SIZE + ECCBITS{1'b0}};
            r[7] = {WORD_SIZE + ECCBITS{1'b0}};
            r[8] = {WORD_SIZE + ECCBITS{1'b0}};
            r[9] = {WORD_SIZE + ECCBITS{1'b0}};
            r[10] = {WORD_SIZE + ECCBITS{1'b0}};
            r[11] = {WORD_SIZE + ECCBITS{1'b0}};
            r[12] = {WORD_SIZE + ECCBITS{1'b0}};
            r[13] = {WORD_SIZE + ECCBITS{1'b0}};
            r[14] = {WORD_SIZE + ECCBITS{1'b0}};
            r[15] = {WORD_SIZE + ECCBITS{1'b0}};
            r[16] = {WORD_SIZE + ECCBITS{1'b0}};
            r[17] = {WORD_SIZE + ECCBITS{1'b0}};
            r[18] = {WORD_SIZE + ECCBITS{1'b0}};
            r[19] = {WORD_SIZE + ECCBITS{1'b0}};
            r[20] = {WORD_SIZE + ECCBITS{1'b0}};
            r[21] = {WORD_SIZE + ECCBITS{1'b0}};
            r[22] = {WORD_SIZE + ECCBITS{1'b0}};
            r[23] = {WORD_SIZE + ECCBITS{1'b0}};
            r[24] = {WORD_SIZE + ECCBITS{1'b0}};
            r[25] = {WORD_SIZE + ECCBITS{1'b0}};
            r[26] = {WORD_SIZE + ECCBITS{1'b0}};
            r[27] = {WORD_SIZE + ECCBITS{1'b0}};
            r[28] = {WORD_SIZE + ECCBITS{1'b0}};
            r[29] = {WORD_SIZE + ECCBITS{1'b0}};
            r[30] = {WORD_SIZE + ECCBITS{1'b0}};
            r[31] = {WORD_SIZE + ECCBITS{1'b0}};
            ready_o <= 1'b0;
            store_data_o = {WORD_SIZE + ECCBITS {1'b0}};
        end
        else if (rregister_i) begin
            store_data_o = r[register_i];
        end
        else if (wregister_i) begin
            // Sore data
            r[register_i] = data_to_register_i;
            store_data_o = {WORD_SIZE + ECCBITS {1'b0}}; 
        end

    end

    always @(posedge clk_i) begin
        if (valid_i) begin
            case (whisbone_addr_i)
                REGISTERDATA: begin
                    ready_o <= 1'b1;
                    if (wbs_we_i) begin
                        if (wstrb_i[0]) r[31][7:0]   <= wdata_i[7:0];
                        if (wstrb_i[1]) r[31][15:8]  <= wdata_i[15:8];
                        if (wstrb_i[2]) r[31][23:16] <= wdata_i[23:16];
                        if (wstrb_i[3]) r[31][31:24] <= wdata_i[31:24];
                    end
                    else begin
                        rdata_o <= {r[31][31:0]};
                    end
                end
                ADDRBASE + 4: begin ready_o <= 1'b1; end
                ADDRBASE + 8: begin ready_o <= 1'b1; end
                ADDRBASE + 16: begin ready_o <= 1'b1; end
                default: ready_o <= 1'b0;
            endcase
        end
    end
        
endmodule
