VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_64_512_sky130
   CLASS BLOCK ;
   SIZE 822.5 BY 334.94 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 0.0 164.26 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.68 0.0 171.06 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  181.56 0.0 181.94 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 0.0 188.06 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.92 0.0 200.3 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 0.0 205.06 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 0.0 211.86 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 0.0 216.62 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.16 0.0 229.54 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  234.6 0.0 234.98 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  240.04 0.0 240.42 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.16 0.0 246.54 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 252.66 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 0.0 258.1 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  263.84 0.0 264.22 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 0.0 270.34 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 0.0 275.1 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  281.52 0.0 281.9 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 0.0 286.66 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 0.0 293.46 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  298.52 0.0 298.9 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 0.0 310.46 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 0.0 316.58 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  321.64 0.0 322.02 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 0.0 328.14 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  333.2 0.0 333.58 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  340.0 0.0 340.38 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.76 0.0 345.14 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  351.56 0.0 351.94 0.38 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  357.0 0.0 357.38 0.38 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  362.44 0.0 362.82 0.38 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  368.56 0.0 368.94 0.38 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  374.68 0.0 375.06 0.38 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  380.12 0.0 380.5 0.38 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  386.24 0.0 386.62 0.38 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  391.68 0.0 392.06 0.38 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  397.8 0.0 398.18 0.38 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  403.92 0.0 404.3 0.38 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  410.04 0.0 410.42 0.38 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  415.48 0.0 415.86 0.38 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  420.92 0.0 421.3 0.38 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  426.36 0.0 426.74 0.38 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  432.48 0.0 432.86 0.38 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  438.6 0.0 438.98 0.38 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 0.0 444.42 0.38 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  450.16 0.0 450.54 0.38 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  455.6 0.0 455.98 0.38 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  461.72 0.0 462.1 0.38 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  468.52 0.0 468.9 0.38 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  473.28 0.0 473.66 0.38 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  479.4 0.0 479.78 0.38 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  484.84 0.0 485.22 0.38 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  490.96 0.0 491.34 0.38 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  497.08 0.0 497.46 0.38 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  502.52 0.0 502.9 0.38 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  509.32 0.0 509.7 0.38 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  514.76 0.0 515.14 0.38 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  520.88 0.0 521.26 0.38 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  526.32 0.0 526.7 0.38 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  532.44 0.0 532.82 0.38 ;
      END
   END din0[63]
   PIN din0[64]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  537.88 0.0 538.26 0.38 ;
      END
   END din0[64]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  106.08 0.0 106.46 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.2 0.0 112.58 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 154.36 0.38 154.74 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.2 0.38 163.58 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 168.64 0.38 169.02 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 177.48 0.38 177.86 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 183.6 0.38 183.98 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 191.08 0.38 191.46 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 197.2 0.38 197.58 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 51.68 0.38 52.06 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 59.84 0.38 60.22 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 53.72 0.38 54.1 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  117.64 0.0 118.02 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 0.0 124.14 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.88 0.0 130.26 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.64 0.0 135.02 0.38 ;
      END
   END wmask0[3]
   PIN wmask0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  141.44 0.0 141.82 0.38 ;
      END
   END wmask0[4]
   PIN wmask0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 0.0 146.58 0.38 ;
      END
   END wmask0[5]
   PIN wmask0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.0 0.0 153.38 0.38 ;
      END
   END wmask0[6]
   PIN wmask0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 0.38 ;
      END
   END wmask0[7]
   PIN spare_wen0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  543.32 0.0 543.7 0.38 ;
      END
   END spare_wen0[0]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.04 0.0 189.42 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 0.0 199.62 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.48 0.0 228.86 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 0.0 247.9 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.08 0.0 259.46 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 0.0 269.66 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.8 0.0 279.18 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  289.0 0.0 289.38 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 0.0 299.58 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  308.04 0.0 308.42 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.92 0.0 319.3 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 0.0 326.1 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  337.28 0.0 337.66 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.84 0.0 349.22 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.04 0.0 359.42 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  369.24 0.0 369.62 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  378.08 0.0 378.46 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  388.96 0.0 389.34 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  399.16 0.0 399.54 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.32 0.0 407.7 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  418.88 0.0 419.26 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  429.08 0.0 429.46 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  439.28 0.0 439.66 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  448.12 0.0 448.5 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  459.0 0.0 459.38 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  469.2 0.0 469.58 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  477.36 0.0 477.74 0.38 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  487.56 0.0 487.94 0.38 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  499.12 0.0 499.5 0.38 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  508.64 0.0 509.02 0.38 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  518.16 0.0 518.54 0.38 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  529.04 0.0 529.42 0.38 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  538.56 0.0 538.94 0.38 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  547.4 0.0 547.78 0.38 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  558.96 0.0 559.34 0.38 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  567.8 0.0 568.18 0.38 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  578.68 0.0 579.06 0.38 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  588.88 0.0 589.26 0.38 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  599.08 0.0 599.46 0.38 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  608.6 0.0 608.98 0.38 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  618.8 0.0 619.18 0.38 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  629.0 0.0 629.38 0.38 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  638.52 0.0 638.9 0.38 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  647.36 0.0 647.74 0.38 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  658.92 0.0 659.3 0.38 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  669.12 0.0 669.5 0.38 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  678.64 0.0 679.02 0.38 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  688.84 0.0 689.22 0.38 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  699.04 0.0 699.42 0.38 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  708.56 0.0 708.94 0.38 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  718.76 0.0 719.14 0.38 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  727.6 0.0 727.98 0.38 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  739.16 0.0 739.54 0.38 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  748.68 0.0 749.06 0.38 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 74.12 822.5 74.5 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 80.24 822.5 80.62 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 79.56 822.5 79.94 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 74.8 822.5 75.18 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 75.48 822.5 75.86 ;
      END
   END dout0[63]
   PIN dout0[64]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  822.12 76.84 822.5 77.22 ;
      END
   END dout0[64]
   PIN vpwr
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 1.36 3.1 334.94 ;
         LAYER met3 ;
         RECT  1.36 1.36 821.14 3.1 ;
         LAYER met4 ;
         RECT  819.4 1.36 821.14 334.94 ;
         LAYER met3 ;
         RECT  1.36 333.2 821.14 334.94 ;
      END
   END vpwr
   PIN vgnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 817.74 6.5 ;
         LAYER met3 ;
         RECT  4.76 329.8 817.74 331.54 ;
         LAYER met4 ;
         RECT  816.0 4.76 817.74 331.54 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 331.54 ;
      END
   END vgnd
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 821.88 334.32 ;
   LAYER  met2 ;
      RECT  0.62 0.62 821.88 334.32 ;
   LAYER  met3 ;
      RECT  0.98 153.76 821.88 155.34 ;
      RECT  0.62 155.34 0.98 162.6 ;
      RECT  0.62 164.18 0.98 168.04 ;
      RECT  0.62 169.62 0.98 176.88 ;
      RECT  0.62 178.46 0.98 183.0 ;
      RECT  0.62 184.58 0.98 190.48 ;
      RECT  0.62 192.06 0.98 196.6 ;
      RECT  0.62 60.82 0.98 153.76 ;
      RECT  0.62 52.66 0.98 53.12 ;
      RECT  0.62 54.7 0.98 59.24 ;
      RECT  0.98 73.52 821.52 75.1 ;
      RECT  0.98 75.1 821.52 153.76 ;
      RECT  821.52 81.22 821.88 153.76 ;
      RECT  821.52 77.82 821.88 78.96 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 51.08 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 51.08 ;
      RECT  0.98 0.62 821.52 0.76 ;
      RECT  821.52 0.62 821.74 0.76 ;
      RECT  821.52 3.7 821.74 73.52 ;
      RECT  821.74 0.62 821.88 0.76 ;
      RECT  821.74 0.76 821.88 3.7 ;
      RECT  821.74 3.7 821.88 73.52 ;
      RECT  821.74 155.34 821.88 332.6 ;
      RECT  821.74 332.6 821.88 334.32 ;
      RECT  0.62 198.18 0.76 332.6 ;
      RECT  0.62 332.6 0.76 334.32 ;
      RECT  0.76 198.18 0.98 332.6 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 73.52 ;
      RECT  4.16 3.7 818.34 4.16 ;
      RECT  4.16 7.1 818.34 73.52 ;
      RECT  818.34 3.7 821.52 4.16 ;
      RECT  818.34 4.16 821.52 7.1 ;
      RECT  818.34 7.1 821.52 73.52 ;
      RECT  0.98 155.34 4.16 329.2 ;
      RECT  0.98 329.2 4.16 332.14 ;
      RECT  0.98 332.14 4.16 332.6 ;
      RECT  4.16 155.34 818.34 329.2 ;
      RECT  4.16 332.14 818.34 332.6 ;
      RECT  818.34 155.34 821.74 329.2 ;
      RECT  818.34 329.2 821.74 332.14 ;
      RECT  818.34 332.14 821.74 332.6 ;
   LAYER  met4 ;
      RECT  163.28 0.98 164.86 334.32 ;
      RECT  171.66 0.62 175.52 0.98 ;
      RECT  182.54 0.62 187.08 0.98 ;
      RECT  200.9 0.62 204.08 0.98 ;
      RECT  212.46 0.62 215.64 0.98 ;
      RECT  230.14 0.62 234.0 0.98 ;
      RECT  241.02 0.62 245.56 0.98 ;
      RECT  253.26 0.62 257.12 0.98 ;
      RECT  270.94 0.62 274.12 0.98 ;
      RECT  282.5 0.62 285.68 0.98 ;
      RECT  294.06 0.62 297.92 0.98 ;
      RECT  311.06 0.62 315.6 0.98 ;
      RECT  328.74 0.62 332.6 0.98 ;
      RECT  340.98 0.62 344.16 0.98 ;
      RECT  352.54 0.62 356.4 0.98 ;
      RECT  363.42 0.62 367.96 0.98 ;
      RECT  381.1 0.62 385.64 0.98 ;
      RECT  392.66 0.62 397.2 0.98 ;
      RECT  411.02 0.62 414.88 0.98 ;
      RECT  421.9 0.62 425.76 0.98 ;
      RECT  433.46 0.62 438.0 0.98 ;
      RECT  451.14 0.62 455.0 0.98 ;
      RECT  462.7 0.62 467.92 0.98 ;
      RECT  480.38 0.62 484.24 0.98 ;
      RECT  491.94 0.62 496.48 0.98 ;
      RECT  510.3 0.62 514.16 0.98 ;
      RECT  521.86 0.62 525.72 0.98 ;
      RECT  533.42 0.62 537.28 0.98 ;
      RECT  107.06 0.62 111.6 0.98 ;
      RECT  113.18 0.62 117.04 0.98 ;
      RECT  118.62 0.62 123.16 0.98 ;
      RECT  124.74 0.62 129.28 0.98 ;
      RECT  130.86 0.62 134.04 0.98 ;
      RECT  135.62 0.62 140.84 0.98 ;
      RECT  142.42 0.62 145.6 0.98 ;
      RECT  147.18 0.62 152.4 0.98 ;
      RECT  153.98 0.62 157.16 0.98 ;
      RECT  158.74 0.62 163.28 0.98 ;
      RECT  164.86 0.62 166.68 0.98 ;
      RECT  168.26 0.62 170.08 0.98 ;
      RECT  177.1 0.62 178.24 0.98 ;
      RECT  179.82 0.62 180.96 0.98 ;
      RECT  190.02 0.62 192.52 0.98 ;
      RECT  194.1 0.62 198.64 0.98 ;
      RECT  205.66 0.62 208.16 0.98 ;
      RECT  209.74 0.62 210.88 0.98 ;
      RECT  217.22 0.62 218.36 0.98 ;
      RECT  219.94 0.62 222.44 0.98 ;
      RECT  224.02 0.62 227.88 0.98 ;
      RECT  235.58 0.62 237.4 0.98 ;
      RECT  238.98 0.62 239.44 0.98 ;
      RECT  248.5 0.62 251.68 0.98 ;
      RECT  260.06 0.62 263.24 0.98 ;
      RECT  264.82 0.62 268.68 0.98 ;
      RECT  275.7 0.62 278.2 0.98 ;
      RECT  279.78 0.62 280.92 0.98 ;
      RECT  287.26 0.62 288.4 0.98 ;
      RECT  289.98 0.62 292.48 0.98 ;
      RECT  300.18 0.62 304.04 0.98 ;
      RECT  305.62 0.62 307.44 0.98 ;
      RECT  309.02 0.62 309.48 0.98 ;
      RECT  317.18 0.62 318.32 0.98 ;
      RECT  319.9 0.62 321.04 0.98 ;
      RECT  322.62 0.62 325.12 0.98 ;
      RECT  326.7 0.62 327.16 0.98 ;
      RECT  334.18 0.62 336.68 0.98 ;
      RECT  338.26 0.62 339.4 0.98 ;
      RECT  345.74 0.62 348.24 0.98 ;
      RECT  349.82 0.62 350.96 0.98 ;
      RECT  357.98 0.62 358.44 0.98 ;
      RECT  360.02 0.62 361.84 0.98 ;
      RECT  370.22 0.62 374.08 0.98 ;
      RECT  375.66 0.62 377.48 0.98 ;
      RECT  379.06 0.62 379.52 0.98 ;
      RECT  387.22 0.62 388.36 0.98 ;
      RECT  389.94 0.62 391.08 0.98 ;
      RECT  400.14 0.62 403.32 0.98 ;
      RECT  404.9 0.62 406.72 0.98 ;
      RECT  408.3 0.62 409.44 0.98 ;
      RECT  416.46 0.62 418.28 0.98 ;
      RECT  419.86 0.62 420.32 0.98 ;
      RECT  427.34 0.62 428.48 0.98 ;
      RECT  430.06 0.62 431.88 0.98 ;
      RECT  440.26 0.62 443.44 0.98 ;
      RECT  445.02 0.62 447.52 0.98 ;
      RECT  449.1 0.62 449.56 0.98 ;
      RECT  456.58 0.62 458.4 0.98 ;
      RECT  459.98 0.62 461.12 0.98 ;
      RECT  470.18 0.62 472.68 0.98 ;
      RECT  474.26 0.62 476.76 0.98 ;
      RECT  478.34 0.62 478.8 0.98 ;
      RECT  485.82 0.62 486.96 0.98 ;
      RECT  488.54 0.62 490.36 0.98 ;
      RECT  498.06 0.62 498.52 0.98 ;
      RECT  500.1 0.62 501.92 0.98 ;
      RECT  503.5 0.62 508.04 0.98 ;
      RECT  515.74 0.62 517.56 0.98 ;
      RECT  519.14 0.62 520.28 0.98 ;
      RECT  527.3 0.62 528.44 0.98 ;
      RECT  530.02 0.62 531.84 0.98 ;
      RECT  539.54 0.62 542.72 0.98 ;
      RECT  544.3 0.62 546.8 0.98 ;
      RECT  548.38 0.62 558.36 0.98 ;
      RECT  559.94 0.62 567.2 0.98 ;
      RECT  568.78 0.62 578.08 0.98 ;
      RECT  579.66 0.62 588.28 0.98 ;
      RECT  589.86 0.62 598.48 0.98 ;
      RECT  600.06 0.62 608.0 0.98 ;
      RECT  609.58 0.62 618.2 0.98 ;
      RECT  619.78 0.62 628.4 0.98 ;
      RECT  629.98 0.62 637.92 0.98 ;
      RECT  639.5 0.62 646.76 0.98 ;
      RECT  648.34 0.62 658.32 0.98 ;
      RECT  659.9 0.62 668.52 0.98 ;
      RECT  670.1 0.62 678.04 0.98 ;
      RECT  679.62 0.62 688.24 0.98 ;
      RECT  689.82 0.62 698.44 0.98 ;
      RECT  700.02 0.62 707.96 0.98 ;
      RECT  709.54 0.62 718.16 0.98 ;
      RECT  719.74 0.62 727.0 0.98 ;
      RECT  728.58 0.62 738.56 0.98 ;
      RECT  740.14 0.62 748.08 0.98 ;
      RECT  0.62 0.98 0.76 334.32 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 105.48 0.76 ;
      RECT  3.7 0.76 105.48 0.98 ;
      RECT  821.74 0.98 821.88 334.32 ;
      RECT  749.66 0.62 818.8 0.76 ;
      RECT  749.66 0.76 818.8 0.98 ;
      RECT  818.8 0.62 821.74 0.76 ;
      RECT  821.74 0.62 821.88 0.76 ;
      RECT  821.74 0.76 821.88 0.98 ;
      RECT  164.86 0.98 815.4 4.16 ;
      RECT  164.86 4.16 815.4 332.14 ;
      RECT  164.86 332.14 815.4 334.32 ;
      RECT  815.4 0.98 818.34 4.16 ;
      RECT  815.4 332.14 818.34 334.32 ;
      RECT  818.34 0.98 818.8 4.16 ;
      RECT  818.34 4.16 818.8 332.14 ;
      RECT  818.34 332.14 818.8 334.32 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 332.14 ;
      RECT  3.7 332.14 4.16 334.32 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 332.14 7.1 334.32 ;
      RECT  7.1 0.98 163.28 4.16 ;
      RECT  7.1 4.16 163.28 332.14 ;
      RECT  7.1 332.14 163.28 334.32 ;
   END
END    sram_1rw0r0w_64_512_sky130
END    LIBRARY
