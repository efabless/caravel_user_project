VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw0r0w_32_1024_sky130
   CLASS BLOCK ;
   SIZE 800.74 BY 347.18 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  124.44 0.0 124.82 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.24 0.0 131.62 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.0 0.0 136.38 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 0.0 142.5 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.92 0.0 149.3 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.68 0.0 154.06 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.48 0.0 160.86 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.24 0.0 165.62 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.04 0.0 172.42 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.16 0.0 178.54 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.6 0.0 183.98 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.72 0.0 190.1 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.16 0.0 195.54 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.28 0.0 201.66 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.04 0.0 206.42 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 0.0 213.22 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.08 0.0 242.46 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 0.0 248.58 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.64 0.0 254.02 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 0.0 260.14 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.52 0.0 264.9 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.32 0.0 271.7 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 0.0 282.58 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.32 0.0 288.7 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.76 0.0 294.14 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 0.0 300.94 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  305.32 0.0 305.7 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  312.12 0.0 312.5 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  83.64 0.0 84.02 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  89.76 0.0 90.14 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  95.2 0.0 95.58 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.96 0.38 168.34 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 175.44 0.38 175.82 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 181.56 0.38 181.94 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 189.72 0.38 190.1 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 196.52 0.38 196.9 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 204.68 0.38 205.06 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 209.44 0.38 209.82 ;
      END
   END addr0[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 64.6 0.38 64.98 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 73.44 0.38 73.82 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 65.28 0.38 65.66 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  101.32 0.0 101.7 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.44 0.0 107.82 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.56 0.0 113.94 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 0.0 120.06 0.38 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 0.0 317.94 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  145.52 0.0 145.9 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.0 0.0 187.38 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 0.0 207.78 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.12 0.0 227.5 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 0.0 247.9 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.24 0.0 267.62 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 0.0 286.66 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.0 0.0 306.38 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  327.08 0.0 327.46 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  346.8 0.0 347.18 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 0.0 367.58 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  386.92 0.0 387.3 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  407.32 0.0 407.7 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  427.04 0.0 427.42 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  446.76 0.0 447.14 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  465.8 0.0 466.18 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  486.88 0.0 487.26 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  507.28 0.0 507.66 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  527.0 0.0 527.38 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  546.72 0.0 547.1 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  567.12 0.0 567.5 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  586.84 0.0 587.22 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  607.24 0.0 607.62 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  625.6 0.0 625.98 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  646.68 0.0 647.06 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  667.08 0.0 667.46 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  686.8 0.0 687.18 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  707.2 0.0 707.58 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  800.36 90.44 800.74 90.82 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  800.36 84.32 800.74 84.7 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  800.36 89.76 800.74 90.14 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  800.36 85.0 800.74 85.38 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 1.36 3.1 347.18 ;
         LAYER met3 ;
         RECT  1.36 1.36 799.38 3.1 ;
         LAYER met4 ;
         RECT  797.64 1.36 799.38 347.18 ;
         LAYER met3 ;
         RECT  1.36 345.44 799.38 347.18 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 795.98 6.5 ;
         LAYER met4 ;
         RECT  794.24 4.76 795.98 343.78 ;
         LAYER met3 ;
         RECT  4.76 342.04 795.98 343.78 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 343.78 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 800.12 346.56 ;
   LAYER  met2 ;
      RECT  0.62 0.62 800.12 346.56 ;
   LAYER  met3 ;
      RECT  0.98 167.36 800.12 168.94 ;
      RECT  0.62 168.94 0.98 174.84 ;
      RECT  0.62 176.42 0.98 180.96 ;
      RECT  0.62 182.54 0.98 189.12 ;
      RECT  0.62 190.7 0.98 195.92 ;
      RECT  0.62 197.5 0.98 204.08 ;
      RECT  0.62 205.66 0.98 208.84 ;
      RECT  0.62 74.42 0.98 167.36 ;
      RECT  0.62 66.26 0.98 72.84 ;
      RECT  0.98 89.84 799.76 91.42 ;
      RECT  0.98 91.42 799.76 167.36 ;
      RECT  799.76 91.42 800.12 167.36 ;
      RECT  799.76 85.98 800.12 89.16 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 64.0 ;
      RECT  0.76 0.62 0.98 0.76 ;
      RECT  0.76 3.7 0.98 64.0 ;
      RECT  0.98 0.62 799.76 0.76 ;
      RECT  799.76 0.62 799.98 0.76 ;
      RECT  799.76 3.7 799.98 83.72 ;
      RECT  799.98 0.62 800.12 0.76 ;
      RECT  799.98 0.76 800.12 3.7 ;
      RECT  799.98 3.7 800.12 83.72 ;
      RECT  799.98 168.94 800.12 344.84 ;
      RECT  799.98 344.84 800.12 346.56 ;
      RECT  0.62 210.42 0.76 344.84 ;
      RECT  0.62 344.84 0.76 346.56 ;
      RECT  0.76 210.42 0.98 344.84 ;
      RECT  0.98 3.7 4.16 4.16 ;
      RECT  0.98 4.16 4.16 7.1 ;
      RECT  0.98 7.1 4.16 89.84 ;
      RECT  4.16 3.7 796.58 4.16 ;
      RECT  4.16 7.1 796.58 89.84 ;
      RECT  796.58 3.7 799.76 4.16 ;
      RECT  796.58 4.16 799.76 7.1 ;
      RECT  796.58 7.1 799.76 89.84 ;
      RECT  0.98 168.94 4.16 341.44 ;
      RECT  0.98 341.44 4.16 344.38 ;
      RECT  0.98 344.38 4.16 344.84 ;
      RECT  4.16 168.94 796.58 341.44 ;
      RECT  4.16 344.38 796.58 344.84 ;
      RECT  796.58 168.94 799.98 341.44 ;
      RECT  796.58 341.44 799.98 344.38 ;
      RECT  796.58 344.38 799.98 344.84 ;
   LAYER  met4 ;
      RECT  123.84 0.98 125.42 346.56 ;
      RECT  125.42 0.62 130.64 0.98 ;
      RECT  132.22 0.62 135.4 0.98 ;
      RECT  136.98 0.62 141.52 0.98 ;
      RECT  149.9 0.62 153.08 0.98 ;
      RECT  154.66 0.62 159.88 0.98 ;
      RECT  161.46 0.62 164.64 0.98 ;
      RECT  173.02 0.62 177.56 0.98 ;
      RECT  179.14 0.62 183.0 0.98 ;
      RECT  190.7 0.62 194.56 0.98 ;
      RECT  196.14 0.62 200.68 0.98 ;
      RECT  202.26 0.62 205.44 0.98 ;
      RECT  213.82 0.62 218.36 0.98 ;
      RECT  219.94 0.62 223.8 0.98 ;
      RECT  231.5 0.62 235.36 0.98 ;
      RECT  236.94 0.62 241.48 0.98 ;
      RECT  249.18 0.62 253.04 0.98 ;
      RECT  254.62 0.62 259.16 0.98 ;
      RECT  260.74 0.62 263.92 0.98 ;
      RECT  272.3 0.62 275.48 0.98 ;
      RECT  277.06 0.62 281.6 0.98 ;
      RECT  289.3 0.62 293.16 0.98 ;
      RECT  294.74 0.62 299.96 0.98 ;
      RECT  301.54 0.62 304.72 0.98 ;
      RECT  84.62 0.62 89.16 0.98 ;
      RECT  90.74 0.62 94.6 0.98 ;
      RECT  96.18 0.62 100.72 0.98 ;
      RECT  102.3 0.62 106.84 0.98 ;
      RECT  108.42 0.62 112.96 0.98 ;
      RECT  114.54 0.62 119.08 0.98 ;
      RECT  120.66 0.62 123.84 0.98 ;
      RECT  313.1 0.62 316.96 0.98 ;
      RECT  143.1 0.62 144.92 0.98 ;
      RECT  146.5 0.62 148.32 0.98 ;
      RECT  166.22 0.62 166.68 0.98 ;
      RECT  168.26 0.62 171.44 0.98 ;
      RECT  184.58 0.62 186.4 0.98 ;
      RECT  187.98 0.62 189.12 0.98 ;
      RECT  208.38 0.62 212.24 0.98 ;
      RECT  225.38 0.62 226.52 0.98 ;
      RECT  228.1 0.62 229.92 0.98 ;
      RECT  243.06 0.62 246.92 0.98 ;
      RECT  265.5 0.62 266.64 0.98 ;
      RECT  268.22 0.62 270.72 0.98 ;
      RECT  283.18 0.62 285.68 0.98 ;
      RECT  287.26 0.62 287.72 0.98 ;
      RECT  306.98 0.62 311.52 0.98 ;
      RECT  318.54 0.62 326.48 0.98 ;
      RECT  328.06 0.62 346.2 0.98 ;
      RECT  347.78 0.62 366.6 0.98 ;
      RECT  368.18 0.62 386.32 0.98 ;
      RECT  387.9 0.62 406.72 0.98 ;
      RECT  408.3 0.62 426.44 0.98 ;
      RECT  428.02 0.62 446.16 0.98 ;
      RECT  447.74 0.62 465.2 0.98 ;
      RECT  466.78 0.62 486.28 0.98 ;
      RECT  487.86 0.62 506.68 0.98 ;
      RECT  508.26 0.62 526.4 0.98 ;
      RECT  527.98 0.62 546.12 0.98 ;
      RECT  547.7 0.62 566.52 0.98 ;
      RECT  568.1 0.62 586.24 0.98 ;
      RECT  587.82 0.62 606.64 0.98 ;
      RECT  608.22 0.62 625.0 0.98 ;
      RECT  626.58 0.62 646.08 0.98 ;
      RECT  647.66 0.62 666.48 0.98 ;
      RECT  668.06 0.62 686.2 0.98 ;
      RECT  687.78 0.62 706.6 0.98 ;
      RECT  0.62 0.98 0.76 346.56 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 0.98 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 83.04 0.76 ;
      RECT  3.7 0.76 83.04 0.98 ;
      RECT  799.98 0.98 800.12 346.56 ;
      RECT  708.18 0.62 797.04 0.76 ;
      RECT  708.18 0.76 797.04 0.98 ;
      RECT  797.04 0.62 799.98 0.76 ;
      RECT  799.98 0.62 800.12 0.76 ;
      RECT  799.98 0.76 800.12 0.98 ;
      RECT  125.42 0.98 793.64 4.16 ;
      RECT  125.42 4.16 793.64 344.38 ;
      RECT  125.42 344.38 793.64 346.56 ;
      RECT  793.64 0.98 796.58 4.16 ;
      RECT  793.64 344.38 796.58 346.56 ;
      RECT  796.58 0.98 797.04 4.16 ;
      RECT  796.58 4.16 797.04 344.38 ;
      RECT  796.58 344.38 797.04 346.56 ;
      RECT  3.7 0.98 4.16 4.16 ;
      RECT  3.7 4.16 4.16 344.38 ;
      RECT  3.7 344.38 4.16 346.56 ;
      RECT  4.16 0.98 7.1 4.16 ;
      RECT  4.16 344.38 7.1 346.56 ;
      RECT  7.1 0.98 123.84 4.16 ;
      RECT  7.1 4.16 123.84 344.38 ;
      RECT  7.1 344.38 123.84 346.56 ;
   END
END    sram_1rw0r0w_32_1024_sky130
END    LIBRARY
