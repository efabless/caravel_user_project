`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***

//***Module***


module register_file #(
        parameter integer WORD_SIZE = 32,
        parameter integer REGISTERS = 32,
        parameter integer REGDIRSIZE = 5,
        parameter integer ECCBITS = 7,
        parameter integer WHISBONE_ADR = 32,
        parameter integer VERIFICATION_PINS = 2,
        parameter integer COUNTERSIZE = 8
    )
    (

        input  clk_i ,
        input  rst_i ,
        // whishbone interface
        input valid_i,
        input [3:0] wstrb_i,
        input [WORD_SIZE - 1 : 0] wdata_i,
        input [WHISBONE_ADR - 1 : 0] whisbone_addr_i,
        input wbs_we_i,
        // end whishbone interface
        input  [WORD_SIZE - 1 : 0] data_to_register_i ,
        input  [REGDIRSIZE - 1 : 0] register_i ,
        input  wregister_i ,
        input  rregister_i ,
        output [WORD_SIZE - 1 : 0] store_data_o ,
        output [VERIFICATION_PINS - 1 : 0] operation_result_o, 
        // whishbone interface
        output ready_o,
        output [WORD_SIZE - 1 : 0] rdata_o
        // end whishbone interface
    );

//***Internal logic generated by compiler***  
    wire [WORD_SIZE + ECCBITS- 1 : 0] data_to_register_PCW_RD; // wiring between data_to_register_o of module PCW and data_to_register_i of module RD
    wire [WORD_SIZE + ECCBITS - 1 : 0] store_data_RD_DV; // wiring between store_data_o of module RD and internal_data_i of module DV
    wire [VERIFICATION_PINS - 1 : 0] operation_result_DV_PMU; // wiring between operation_result_o of module DV and operation_result_i of module PMU
    wire valid_output_DV_PMU; // wiring between valid_output_o of module DV and valid_output_i of module PMU
    wire [WORD_SIZE - 1 : 0] store_data_DV_DO; // wiring between store_data_o of module DV and store_data_i of module DO

    parity_calculator #(
        .WORD_SIZE (WORD_SIZE),
        .ECCBITS (ECCBITS)
    )
    inst_PCW(
        .data_to_register_i       (data_to_register_i ),
        .operate_i                (wregister_i ),
        .data_to_register_o       (data_to_register_PCW_RD)
    );

    register_data #(
        .WORD_SIZE (WORD_SIZE),
        .REGISTERS (REGISTERS),
        .REGDIRSIZE (REGDIRSIZE),
        .ECCBITS (ECCBITS),
        .WHISBONE_ADR (WHISBONE_ADR)

    )
    inst_RD(
        .clk_i                     (clk_i ),
        .rst_i                     (rst_i ),
        .data_to_register_i        (data_to_register_PCW_RD),
        .register_i                (register_i ),
        .wregister_i               (wregister_i ),
        .rregister_i               (rregister_i ),
        .valid_i                   (valid_i),
        .wstrb_i                   (wstrb_i),
        .wbs_we_i                  (wbs_we_i),
        .wdata_i                   (wdata_i),
        .whisbone_addr_i           (whisbone_addr_i),
        .store_data_o              (store_data_RD_DV),
        .ready_o                   (ready_o),
        .rdata_o                   (rdata_o)
    );

    data_verificator #(
        .WORD_SIZE (WORD_SIZE),
        .ECCBITS (ECCBITS),
        .VERIFICATION_PINS (VERIFICATION_PINS)
    )
    inst_DV(
        .internal_data_i          (store_data_RD_DV),
        .operate_i                (rregister_i ),
        .operation_result_o       (operation_result_DV_PMU),
        .store_data_o             (store_data_DV_DO),
        .valid_output_o           (valid_output_DV_PMU)
    );

    decoder_output #(
        .WORD_SIZE (WORD_SIZE)
    )
    inst_DO(
        .operation_result_i       (operation_result_DV_PMU),
        .store_data_i             (store_data_DV_DO),
        .operation_result_o       (operation_result_o ),
        .store_data_o             (store_data_o )
    );

    state_counters #(
        .WORD_SIZE (WORD_SIZE),
        .VERIFICATION_PINS (VERIFICATION_PINS),
        .WHISBONE_ADR (WHISBONE_ADR),
        .COUNTERSIZE (COUNTERSIZE)
    )
    inst_PMU(
        .clk_i                    (clk_i ),
        .rst_i                    (rst_i ),
        .valid_i                  (valid_i),
        .wstrb_i                  (wstrb_i),
        .wdata_i                  (wdata_i),
        .wbs_we_i                 (wbs_we_i),
        .whisbone_addr_i          (whisbone_addr_i),
        .operation_result_i       (operation_result_DV_PMU),
        .valid_output_i           (valid_output_DV_PMU),
        .ready_o                  (ready_o),
        .rdata_o                  (rdata_o)
    );


//***Handcrafted Internal logic*** 
//TODO
endmodule
