* SPICE3 file created from /home/sky/asyn_rst_8_gray_counter.ext - technology: sky130A

.option scale=5000u

.subckt x/home/sky/asyn_rst_8_gray_counter RSTB CLK Vdd gnd
C0 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# 2.74fF
C1 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# 2.74fF
C2 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# 2.74fF
C3 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# 2.74fF
C4 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# 2.74fF
C5 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# 2.74fF
C6 Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B 2.66fF
C7 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# 2.74fF
C8 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# 2.74fF
C9 Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B 2.67fF
C10 asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B Vdd 2.67fF
C11 asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B Vdd 2.04fF
C12 Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B 2.67fF
C13 Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B 2.29fF
C14 asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B Vdd 2.67fF
C15 asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B Vdd 2.66fF
C16 CLK RSTB 11.73fF
C17 Vdd RSTB 14.13fF
Xasyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
XT_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B sky130_fd_sc_lp__dfrtp_1
XT_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A
+ T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
XT_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A
+ T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
XT_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A
+ T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
XT_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A
+ T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
XT_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B sky130_fd_sc_lp__dfrtp_1
XT_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B sky130_fd_sc_lp__dfrtp_1
XT_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0 asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B
+ sky130_fd_sc_lp__and2_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3 CLK asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_0 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_1 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_2 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B
+ asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd gnd Vdd Vdd asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ sky130_fd_sc_lp__xor2_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_0 CLK asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_1 CLK asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
Xasyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_2 CLK asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/X
+ RSTB gnd gnd Vdd Vdd asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B sky130_fd_sc_lp__dfrtp_1
C18 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C19 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C20 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C21 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C22 asyn_rst_counter_cell_0/sky130_fd_sc_lp__and2_1_0/B gnd 2.55fF
C23 asyn_rst_counter_cell_0/sky130_fd_sc_lp__xor2_1_0/B gnd 7.64fF
C24 asyn_rst_counter_cell_0/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C25 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.16fF **FLOATING
C26 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C27 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C28 T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C29 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/A gnd 2.91fF
C30 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/B gnd 5.51fF
C31 T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.01fF **FLOATING
C32 CLK gnd 17.70fF
C33 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.16fF **FLOATING
C34 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C35 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C36 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C37 Vdd gnd 177.13fF
C38 asyn_rst_counter_cell_6/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C39 asyn_rst_counter_cell_6/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C40 asyn_rst_counter_cell_6/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C41 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C42 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C43 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C44 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C45 asyn_rst_counter_cell_5/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C46 asyn_rst_counter_cell_5/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C47 asyn_rst_counter_cell_5/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C48 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C49 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C50 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C51 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C52 asyn_rst_counter_cell_4/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C53 asyn_rst_counter_cell_4/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C54 asyn_rst_counter_cell_4/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C55 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C56 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C57 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C58 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C59 asyn_rst_counter_cell_3/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C60 asyn_rst_counter_cell_3/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C61 asyn_rst_counter_cell_3/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C62 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C63 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C64 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C65 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C66 asyn_rst_counter_cell_2/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C67 asyn_rst_counter_cell_2/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C68 asyn_rst_counter_cell_2/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
C69 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_559_533# gnd 2.26fF **FLOATING
C70 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_695_375# gnd 2.62fF **FLOATING
C71 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_27_114# gnd 7.42fF **FLOATING
C72 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__dfrtp_1_3/a_196_462# gnd 4.48fF **FLOATING
C73 asyn_rst_counter_cell_1/sky130_fd_sc_lp__and2_1_0/B gnd 3.25fF
C74 asyn_rst_counter_cell_1/sky130_fd_sc_lp__xor2_1_0/B gnd 8.70fF
C75 asyn_rst_counter_cell_1/T_flip_flop_0/sky130_fd_sc_lp__xor2_1_3/a_42_367# gnd 3.03fF **FLOATING
.ends
