magic
tech sky130A
magscale 1 2
timestamp 1640851109
<< pwell >>
rect 8093 120 8177 234
<< ndiff >>
rect 8142 156 8151 172
<< poly >>
rect 71 265 87 333
rect 842 292 882 337
<< locali >>
rect 23 408 73 415
rect 23 374 34 408
rect 68 374 73 408
rect 23 363 73 374
rect 24 313 74 320
rect 24 279 35 313
rect 69 279 74 313
rect 24 268 74 279
rect 1204 260 1238 272
<< viali >>
rect 2726 491 2760 531
rect 4358 487 4392 521
rect 8762 502 8804 541
rect 34 374 68 408
rect 188 359 222 394
rect 940 350 974 384
rect 5989 357 6026 391
rect 35 279 69 313
rect 392 311 426 345
rect 648 294 682 328
rect 842 292 882 337
rect 1202 272 1240 308
rect 1521 269 1563 316
rect 3143 274 3183 320
rect 2840 202 2876 241
rect 4459 240 4498 279
rect 4779 275 4819 318
rect 6412 279 6450 321
rect 6089 240 6126 279
rect 7739 277 7779 312
rect 8386 298 8439 359
rect 8576 346 8621 395
rect 7908 242 7943 277
rect 7621 136 7656 171
rect 8117 156 8151 191
<< metal1 >>
rect 176 564 1132 592
rect 176 528 208 564
rect 0 496 208 528
rect 18 417 86 428
rect 18 404 24 417
rect 0 372 24 404
rect 18 365 24 372
rect 76 365 86 417
rect 176 412 208 496
rect 382 506 1062 534
rect 18 360 86 365
rect 175 394 239 412
rect 175 359 188 394
rect 222 359 239 394
rect 382 362 412 506
rect 930 395 991 407
rect 175 343 239 359
rect 381 345 433 362
rect 19 322 87 332
rect 19 311 25 322
rect 0 279 25 311
rect 19 270 25 279
rect 77 270 87 322
rect 381 311 392 345
rect 426 311 433 345
rect 834 340 893 351
rect 632 330 712 339
rect 381 295 433 311
rect 484 328 712 330
rect 19 265 87 270
rect 484 294 648 328
rect 682 294 712 328
rect 484 284 712 294
rect 484 208 513 284
rect 632 283 712 284
rect 0 176 513 208
rect 680 118 712 283
rect 834 285 838 340
rect 890 285 893 340
rect 930 343 934 395
rect 986 343 991 395
rect 930 331 991 343
rect 834 273 893 285
rect 1020 219 1062 506
rect 1098 326 1132 564
rect 2712 544 2775 554
rect 2712 531 3209 544
rect 2712 491 2726 531
rect 2760 512 3209 531
rect 2760 491 2775 512
rect 2712 447 2775 491
rect 1098 308 1248 326
rect 1098 296 1202 308
rect 1189 272 1202 296
rect 1240 296 1248 308
rect 1500 316 1586 359
rect 1240 272 1247 296
rect 1189 248 1247 272
rect 1500 269 1521 316
rect 1563 269 1586 316
rect 1500 219 1586 269
rect 3120 320 3209 512
rect 4347 525 4410 567
rect 8744 552 8822 582
rect 8744 541 8893 552
rect 4347 521 7798 525
rect 4347 487 4358 521
rect 4392 493 7798 521
rect 4392 487 4410 493
rect 4347 426 4410 487
rect 3120 274 3143 320
rect 3183 274 3209 320
rect 1020 186 1586 219
rect 2818 241 2891 250
rect 2818 202 2840 241
rect 2876 202 2891 241
rect 3120 240 3209 274
rect 4446 279 4512 328
rect 4446 240 4459 279
rect 4498 240 4512 279
rect 2818 118 2891 202
rect 680 117 2891 118
rect 4446 117 4512 240
rect 4750 318 4837 493
rect 7729 440 7798 493
rect 8744 502 8762 541
rect 8804 520 8893 541
rect 8804 502 8822 520
rect 8744 470 8822 502
rect 7729 438 8632 440
rect 5982 391 6040 430
rect 5982 357 5989 391
rect 6026 377 6040 391
rect 7729 428 8639 438
rect 7729 408 8893 428
rect 6026 357 6477 377
rect 5982 330 6477 357
rect 5982 324 6040 330
rect 4750 275 4779 318
rect 4819 275 4837 318
rect 6380 321 6477 330
rect 4750 239 4837 275
rect 6075 279 6149 293
rect 6075 240 6089 279
rect 6126 240 6149 279
rect 6380 279 6412 321
rect 6450 279 6477 321
rect 6380 241 6477 279
rect 7729 312 7798 408
rect 8566 396 8893 408
rect 8566 395 8639 396
rect 7729 277 7739 312
rect 7779 277 7798 312
rect 8378 359 8471 379
rect 6075 117 6149 240
rect 7729 235 7798 277
rect 7864 277 7962 306
rect 7864 242 7908 277
rect 7943 242 7962 277
rect 680 85 6149 117
rect 7610 184 7672 230
rect 7864 184 7962 242
rect 8378 298 8386 359
rect 8439 298 8471 359
rect 8566 346 8576 395
rect 8621 346 8639 395
rect 8566 306 8639 346
rect 7610 171 7962 184
rect 7610 136 7621 171
rect 7656 152 7962 171
rect 7656 136 7672 152
rect 7864 151 7962 152
rect 8093 191 8177 234
rect 8378 233 8471 298
rect 8093 156 8117 191
rect 8151 156 8177 191
rect 7610 93 7672 136
rect 8093 126 8177 156
rect 8385 218 8471 233
rect 8385 186 8893 218
rect 8385 137 8443 186
rect 8385 126 8442 137
rect 8093 94 8442 126
rect 680 84 712 85
rect 6075 84 6149 85
<< via1 >>
rect 24 408 76 417
rect 24 374 34 408
rect 34 374 68 408
rect 68 374 76 408
rect 24 365 76 374
rect 25 313 77 322
rect 25 279 35 313
rect 35 279 69 313
rect 69 279 77 313
rect 25 270 77 279
rect 838 337 890 340
rect 838 292 842 337
rect 842 292 882 337
rect 882 292 890 337
rect 838 285 890 292
rect 934 384 986 395
rect 934 350 940 384
rect 940 350 974 384
rect 974 350 986 384
rect 934 343 986 350
<< metal2 >>
rect 18 417 86 428
rect 18 365 24 417
rect 76 410 86 417
rect 76 395 991 410
rect 76 374 934 395
rect 76 365 86 374
rect 18 360 86 365
rect 833 340 893 346
rect 19 323 87 332
rect 833 323 838 340
rect 19 322 838 323
rect 19 270 25 322
rect 77 287 838 322
rect 77 270 87 287
rect 833 285 838 287
rect 890 285 893 340
rect 929 343 934 374
rect 986 343 991 395
rect 929 332 991 343
rect 833 273 893 285
rect 19 265 87 270
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640850677
transform 1 0 7690 0 1 0
box -38 -49 710 715
use comparator_42_18  comparator_42_18_0
timestamp 1640845691
transform 1 0 186 0 1 282
box -186 -282 976 388
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640415294
transform 1 0 1162 0 1 0
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_1
timestamp 1640415294
transform 1 0 2794 0 1 0
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_2
timestamp 1640415294
transform 1 0 4426 0 1 0
box -38 -49 1670 715
use sky130_fd_sc_lp__dfxtp_1  sky130_fd_sc_lp__dfxtp_1_3
timestamp 1640415294
transform 1 0 6058 0 1 0
box -38 -49 1670 715
use sky130_fd_sc_lp__and2_0  sky130_fd_sc_lp__and2_0_0 ~/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 8362 0 1 0
box -38 -49 518 715
<< labels >>
rlabel metal1 8893 537 8893 537 3 polxevent
rlabel metal1 8893 410 8893 410 3 polarity
rlabel metal1 8893 200 8893 200 3 events
<< end >>
