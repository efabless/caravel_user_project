`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***
//***Module***
module decoder_output #(
        parameter integer WORD_SIZE = 32
    )
    (
        input  clk_i ,
        input  [1 : 0] operation_result_i ,
        input  [WORD_SIZE - 1 : 0] store_data_i ,
        output reg [1 : 0] operation_result_o ,
        output reg [WORD_SIZE - 1 : 0] store_data_o 
    );

//***Internal logic generated by compiler***  
    

//***Dumped Internal logic***
    always @(posedge clk_i) begin
        operation_result_o <= operation_result_i;
        store_data_o <= store_data_i;
    end

    
//***Handcrafted Internal logic*** 
//TODO
endmodule
