magic
tech sky130A
timestamp 1640997824
<< nwell >>
rect 27 121 272 205
<< nmos >>
rect 211 44 226 86
<< pmos >>
rect 211 139 226 181
<< ndiff >>
rect 183 73 211 86
rect 183 56 188 73
rect 205 56 211 73
rect 183 44 211 56
rect 226 73 254 86
rect 226 56 232 73
rect 249 56 254 73
rect 226 44 254 56
<< pdiff >>
rect 183 169 211 181
rect 183 152 188 169
rect 205 152 211 169
rect 183 139 211 152
rect 226 169 254 181
rect 226 152 232 169
rect 249 152 254 169
rect 226 139 254 152
<< ndiffc >>
rect 188 56 205 73
rect 232 56 249 73
<< pdiffc >>
rect 188 152 205 169
rect 232 152 249 169
<< poly >>
rect 199 227 238 232
rect 199 210 209 227
rect 228 210 238 227
rect 199 189 238 210
rect 211 181 226 189
rect 211 86 226 139
rect 211 36 226 44
rect 199 22 238 36
rect 199 5 209 22
rect 228 5 238 22
rect 199 0 238 5
<< polycont >>
rect 209 210 228 227
rect 209 5 228 22
<< locali >>
rect 112 231 132 253
rect 199 231 238 232
rect 112 227 238 231
rect 112 211 209 227
rect 112 120 132 211
rect 199 210 209 211
rect 228 210 238 227
rect 199 198 238 210
rect 183 171 209 181
rect 161 169 209 171
rect 161 152 188 169
rect 205 152 209 169
rect 183 139 209 152
rect 228 169 254 181
rect 228 152 232 169
rect 249 152 254 169
rect 228 139 254 152
rect 84 100 132 120
rect 234 120 254 139
rect 234 100 265 120
rect 234 86 254 100
rect 183 73 209 86
rect 163 56 188 73
rect 205 56 209 73
rect 163 54 209 56
rect 183 44 209 54
rect 228 73 254 86
rect 228 56 232 73
rect 249 56 254 73
rect 228 44 254 56
rect 199 22 238 27
rect 199 5 209 22
rect 228 5 238 22
rect 199 0 238 5
<< viali >>
rect 48 210 67 227
rect 27 152 44 169
rect 188 152 205 169
rect 27 56 44 73
rect 188 56 205 73
rect 48 5 67 22
<< metal1 >>
rect 38 227 77 236
rect 38 210 48 227
rect 67 210 77 227
rect 38 205 77 210
rect 22 171 50 176
rect 183 171 211 177
rect -14 169 211 171
rect -14 152 27 169
rect 44 152 188 169
rect 205 152 211 169
rect 22 145 50 152
rect 183 146 211 152
rect 22 73 50 79
rect 183 73 211 79
rect -13 56 27 73
rect 44 56 188 73
rect 205 56 212 73
rect -13 54 212 56
rect 22 48 50 54
rect 183 48 211 54
rect 38 22 77 27
rect 38 5 48 22
rect 67 5 77 22
rect 38 -3 77 5
use inv_lp  inv_lp_0
timestamp 1640995782
transform 1 0 61 0 1 42
box -61 -42 50 190
<< end >>
