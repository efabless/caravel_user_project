VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_4kbyte_1rw1r_32x1024_8
   CLASS BLOCK ;
   SIZE 693.98 BY 668.82 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.32 0.0 118.7 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.76 0.0 124.14 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.88 0.0 130.26 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  135.32 0.0 135.7 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.76 0.0 141.14 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 0.0 146.58 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.0 0.0 153.38 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.12 0.0 159.5 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  164.56 0.0 164.94 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 0.0 170.38 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  175.44 0.0 175.82 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 0.0 182.62 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 0.0 188.06 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.92 0.0 200.3 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.04 0.0 206.42 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 0.0 211.86 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 0.0 217.3 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  222.36 0.0 222.74 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.16 0.0 229.54 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  234.6 0.0 234.98 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  240.72 0.0 241.1 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.16 0.0 246.54 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  251.6 0.0 251.98 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  258.4 0.0 258.78 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  263.84 0.0 264.22 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 0.0 269.66 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 0.0 275.1 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  281.52 0.0 281.9 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 0.0 288.02 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 0.0 293.46 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  298.52 0.0 298.9 1.06 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.96 0.0 83.34 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.4 0.0 88.78 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.92 1.06 149.3 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.08 1.06 157.46 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.88 1.06 164.26 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 171.36 1.06 171.74 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 176.8 1.06 177.18 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 185.64 1.06 186.02 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 191.08 1.06 191.46 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 200.6 1.06 200.98 ;
      END
   END addr0[9]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  605.88 667.76 606.26 668.82 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  599.76 667.76 600.14 668.82 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  692.92 96.56 693.98 96.94 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  692.92 87.04 693.98 87.42 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  692.92 82.28 693.98 82.66 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  692.92 73.44 693.98 73.82 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  624.24 0.0 624.62 1.06 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  622.2 0.0 622.58 1.06 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  622.88 0.0 623.26 1.06 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  623.56 0.0 623.94 1.06 ;
      END
   END addr1[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 1.06 40.5 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  692.92 649.4 693.98 649.78 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 48.96 1.06 49.34 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 41.48 1.06 41.86 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  663.68 667.76 664.06 668.82 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.84 0.0 94.22 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  100.64 0.0 101.02 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.4 0.0 105.78 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  111.52 0.0 111.9 1.06 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 0.0 145.22 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 0.0 160.18 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.04 0.0 172.42 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.2 0.0 197.58 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.0 0.0 221.38 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  249.56 0.0 249.94 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 0.0 260.14 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 0.0 285.3 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  296.48 0.0 296.86 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.32 0.0 322.7 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.56 0.0 334.94 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  347.48 0.0 347.86 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.72 0.0 360.1 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 0.0 372.34 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  384.2 0.0 384.58 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  397.12 0.0 397.5 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  409.36 0.0 409.74 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  421.6 0.0 421.98 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  434.52 0.0 434.9 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  445.4 0.0 445.78 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  459.68 0.0 460.06 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  471.92 0.0 472.3 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  484.16 0.0 484.54 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  497.08 0.0 497.46 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  509.32 0.0 509.7 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  521.56 0.0 521.94 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  534.48 0.0 534.86 1.06 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 667.76 148.62 668.82 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.8 667.76 160.18 668.82 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 667.76 173.1 668.82 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 667.76 185.34 668.82 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 667.76 198.26 668.82 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 667.76 210.5 668.82 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 667.76 223.42 668.82 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 667.76 235.66 668.82 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.52 667.76 247.9 668.82 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.76 667.76 260.14 668.82 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.0 667.76 272.38 668.82 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.92 667.76 285.3 668.82 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 667.76 298.22 668.82 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 667.76 310.46 668.82 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 667.76 323.38 668.82 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.24 667.76 335.62 668.82 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  346.8 667.76 347.18 668.82 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  360.4 667.76 360.78 668.82 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  371.96 667.76 372.34 668.82 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  384.88 667.76 385.26 668.82 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  397.12 667.76 397.5 668.82 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  410.04 667.76 410.42 668.82 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  422.28 667.76 422.66 668.82 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  435.2 667.76 435.58 668.82 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  447.44 667.76 447.82 668.82 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  459.68 667.76 460.06 668.82 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  471.92 667.76 472.3 668.82 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  484.16 667.76 484.54 668.82 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  497.08 667.76 497.46 668.82 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  510.0 667.76 510.38 668.82 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  522.24 667.76 522.62 668.82 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  535.16 667.76 535.54 668.82 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  4.76 4.76 6.5 664.06 ;
         LAYER met3 ;
         RECT  4.76 4.76 689.22 6.5 ;
         LAYER met4 ;
         RECT  687.48 4.76 689.22 664.06 ;
         LAYER met3 ;
         RECT  4.76 662.32 689.22 664.06 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 1.36 3.1 667.46 ;
         LAYER met3 ;
         RECT  1.36 665.72 692.62 667.46 ;
         LAYER met3 ;
         RECT  1.36 1.36 692.62 3.1 ;
         LAYER met4 ;
         RECT  690.88 1.36 692.62 667.46 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 693.36 668.2 ;
   LAYER  met2 ;
      RECT  0.62 0.62 693.36 668.2 ;
   LAYER  met3 ;
      RECT  1.66 148.32 693.36 149.9 ;
      RECT  0.62 149.9 1.66 156.48 ;
      RECT  0.62 158.06 1.66 163.28 ;
      RECT  0.62 164.86 1.66 170.76 ;
      RECT  0.62 172.34 1.66 176.2 ;
      RECT  0.62 177.78 1.66 185.04 ;
      RECT  0.62 186.62 1.66 190.48 ;
      RECT  0.62 192.06 1.66 200.0 ;
      RECT  1.66 95.96 692.32 97.54 ;
      RECT  1.66 97.54 692.32 148.32 ;
      RECT  692.32 97.54 693.36 148.32 ;
      RECT  692.32 88.02 693.36 95.96 ;
      RECT  692.32 83.26 693.36 86.44 ;
      RECT  692.32 74.42 693.36 81.68 ;
      RECT  1.66 149.9 692.32 648.8 ;
      RECT  1.66 648.8 692.32 650.38 ;
      RECT  692.32 149.9 693.36 648.8 ;
      RECT  0.62 49.94 1.66 148.32 ;
      RECT  0.62 42.46 1.66 48.36 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 95.96 ;
      RECT  4.16 7.1 689.82 95.96 ;
      RECT  689.82 4.16 692.32 7.1 ;
      RECT  689.82 7.1 692.32 95.96 ;
      RECT  1.66 650.38 4.16 661.72 ;
      RECT  1.66 661.72 4.16 664.66 ;
      RECT  4.16 650.38 689.82 661.72 ;
      RECT  689.82 650.38 692.32 661.72 ;
      RECT  689.82 661.72 692.32 664.66 ;
      RECT  0.62 201.58 0.76 665.12 ;
      RECT  0.62 665.12 0.76 668.06 ;
      RECT  0.62 668.06 0.76 668.2 ;
      RECT  0.76 201.58 1.66 665.12 ;
      RECT  0.76 668.06 1.66 668.2 ;
      RECT  692.32 650.38 693.22 665.12 ;
      RECT  692.32 668.06 693.22 668.2 ;
      RECT  693.22 650.38 693.36 665.12 ;
      RECT  693.22 665.12 693.36 668.06 ;
      RECT  693.22 668.06 693.36 668.2 ;
      RECT  1.66 664.66 4.16 665.12 ;
      RECT  1.66 668.06 4.16 668.2 ;
      RECT  4.16 664.66 689.82 665.12 ;
      RECT  4.16 668.06 689.82 668.2 ;
      RECT  689.82 664.66 692.32 665.12 ;
      RECT  689.82 668.06 692.32 668.2 ;
      RECT  692.32 0.62 693.22 0.76 ;
      RECT  692.32 3.7 693.22 72.84 ;
      RECT  693.22 0.62 693.36 0.76 ;
      RECT  693.22 0.76 693.36 3.7 ;
      RECT  693.22 3.7 693.36 72.84 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 39.52 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 39.52 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 689.82 0.76 ;
      RECT  4.16 3.7 689.82 4.16 ;
      RECT  689.82 0.62 692.32 0.76 ;
      RECT  689.82 3.7 692.32 4.16 ;
   LAYER  met4 ;
      RECT  117.72 1.66 119.3 668.2 ;
      RECT  119.3 0.62 123.16 1.66 ;
      RECT  124.74 0.62 129.28 1.66 ;
      RECT  130.86 0.62 134.72 1.66 ;
      RECT  136.3 0.62 140.16 1.66 ;
      RECT  147.18 0.62 152.4 1.66 ;
      RECT  153.98 0.62 158.52 1.66 ;
      RECT  165.54 0.62 169.4 1.66 ;
      RECT  176.42 0.62 181.64 1.66 ;
      RECT  188.66 0.62 192.52 1.66 ;
      RECT  200.9 0.62 205.44 1.66 ;
      RECT  212.46 0.62 216.32 1.66 ;
      RECT  223.34 0.62 228.56 1.66 ;
      RECT  235.58 0.62 240.12 1.66 ;
      RECT  241.7 0.62 245.56 1.66 ;
      RECT  252.58 0.62 257.8 1.66 ;
      RECT  264.82 0.62 268.68 1.66 ;
      RECT  275.7 0.62 280.92 1.66 ;
      RECT  288.62 0.62 292.48 1.66 ;
      RECT  83.94 0.62 87.8 1.66 ;
      RECT  119.3 1.66 605.28 667.16 ;
      RECT  605.28 1.66 606.86 667.16 ;
      RECT  600.74 667.16 605.28 668.2 ;
      RECT  606.86 667.16 663.08 668.2 ;
      RECT  89.38 0.62 93.24 1.66 ;
      RECT  94.82 0.62 100.04 1.66 ;
      RECT  101.62 0.62 104.8 1.66 ;
      RECT  106.38 0.62 110.92 1.66 ;
      RECT  112.5 0.62 117.72 1.66 ;
      RECT  141.74 0.62 144.24 1.66 ;
      RECT  160.78 0.62 163.96 1.66 ;
      RECT  170.98 0.62 171.44 1.66 ;
      RECT  173.02 0.62 174.84 1.66 ;
      RECT  183.22 0.62 184.36 1.66 ;
      RECT  185.94 0.62 187.08 1.66 ;
      RECT  194.1 0.62 196.6 1.66 ;
      RECT  198.18 0.62 199.32 1.66 ;
      RECT  207.02 0.62 208.16 1.66 ;
      RECT  209.74 0.62 210.88 1.66 ;
      RECT  217.9 0.62 220.4 1.66 ;
      RECT  230.14 0.62 231.96 1.66 ;
      RECT  233.54 0.62 234.0 1.66 ;
      RECT  247.14 0.62 248.96 1.66 ;
      RECT  250.54 0.62 251.0 1.66 ;
      RECT  260.74 0.62 263.24 1.66 ;
      RECT  270.26 0.62 272.08 1.66 ;
      RECT  273.66 0.62 274.12 1.66 ;
      RECT  282.5 0.62 284.32 1.66 ;
      RECT  285.9 0.62 287.04 1.66 ;
      RECT  294.06 0.62 295.88 1.66 ;
      RECT  297.46 0.62 297.92 1.66 ;
      RECT  299.5 0.62 308.8 1.66 ;
      RECT  310.38 0.62 321.72 1.66 ;
      RECT  323.3 0.62 333.96 1.66 ;
      RECT  335.54 0.62 346.88 1.66 ;
      RECT  348.46 0.62 359.12 1.66 ;
      RECT  360.7 0.62 371.36 1.66 ;
      RECT  372.94 0.62 383.6 1.66 ;
      RECT  385.18 0.62 396.52 1.66 ;
      RECT  398.1 0.62 408.76 1.66 ;
      RECT  410.34 0.62 421.0 1.66 ;
      RECT  422.58 0.62 433.92 1.66 ;
      RECT  435.5 0.62 444.8 1.66 ;
      RECT  446.38 0.62 459.08 1.66 ;
      RECT  460.66 0.62 471.32 1.66 ;
      RECT  472.9 0.62 483.56 1.66 ;
      RECT  485.14 0.62 496.48 1.66 ;
      RECT  498.06 0.62 508.72 1.66 ;
      RECT  510.3 0.62 520.96 1.66 ;
      RECT  522.54 0.62 533.88 1.66 ;
      RECT  535.46 0.62 621.6 1.66 ;
      RECT  119.3 667.16 147.64 668.2 ;
      RECT  149.22 667.16 159.2 668.2 ;
      RECT  160.78 667.16 172.12 668.2 ;
      RECT  173.7 667.16 184.36 668.2 ;
      RECT  185.94 667.16 197.28 668.2 ;
      RECT  198.86 667.16 209.52 668.2 ;
      RECT  211.1 667.16 222.44 668.2 ;
      RECT  224.02 667.16 234.68 668.2 ;
      RECT  236.26 667.16 246.92 668.2 ;
      RECT  248.5 667.16 259.16 668.2 ;
      RECT  260.74 667.16 271.4 668.2 ;
      RECT  272.98 667.16 284.32 668.2 ;
      RECT  285.9 667.16 297.24 668.2 ;
      RECT  298.82 667.16 309.48 668.2 ;
      RECT  311.06 667.16 322.4 668.2 ;
      RECT  323.98 667.16 334.64 668.2 ;
      RECT  336.22 667.16 346.2 668.2 ;
      RECT  347.78 667.16 359.8 668.2 ;
      RECT  361.38 667.16 371.36 668.2 ;
      RECT  372.94 667.16 384.28 668.2 ;
      RECT  385.86 667.16 396.52 668.2 ;
      RECT  398.1 667.16 409.44 668.2 ;
      RECT  411.02 667.16 421.68 668.2 ;
      RECT  423.26 667.16 434.6 668.2 ;
      RECT  436.18 667.16 446.84 668.2 ;
      RECT  448.42 667.16 459.08 668.2 ;
      RECT  460.66 667.16 471.32 668.2 ;
      RECT  472.9 667.16 483.56 668.2 ;
      RECT  485.14 667.16 496.48 668.2 ;
      RECT  498.06 667.16 509.4 668.2 ;
      RECT  510.98 667.16 521.64 668.2 ;
      RECT  523.22 667.16 534.56 668.2 ;
      RECT  536.14 667.16 599.16 668.2 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 664.66 7.1 668.2 ;
      RECT  7.1 1.66 117.72 4.16 ;
      RECT  7.1 4.16 117.72 664.66 ;
      RECT  7.1 664.66 117.72 668.2 ;
      RECT  606.86 1.66 686.88 4.16 ;
      RECT  606.86 4.16 686.88 664.66 ;
      RECT  606.86 664.66 686.88 667.16 ;
      RECT  686.88 1.66 689.82 4.16 ;
      RECT  686.88 664.66 689.82 667.16 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 82.36 0.76 ;
      RECT  3.7 0.76 82.36 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 664.66 ;
      RECT  3.7 4.16 4.16 664.66 ;
      RECT  0.62 664.66 0.76 668.06 ;
      RECT  0.62 668.06 0.76 668.2 ;
      RECT  0.76 668.06 3.7 668.2 ;
      RECT  3.7 664.66 4.16 668.06 ;
      RECT  3.7 668.06 4.16 668.2 ;
      RECT  625.22 0.62 690.28 0.76 ;
      RECT  625.22 0.76 690.28 1.66 ;
      RECT  690.28 0.62 693.22 0.76 ;
      RECT  693.22 0.62 693.36 0.76 ;
      RECT  693.22 0.76 693.36 1.66 ;
      RECT  664.66 667.16 690.28 668.06 ;
      RECT  664.66 668.06 690.28 668.2 ;
      RECT  690.28 668.06 693.22 668.2 ;
      RECT  693.22 667.16 693.36 668.06 ;
      RECT  693.22 668.06 693.36 668.2 ;
      RECT  689.82 1.66 690.28 4.16 ;
      RECT  693.22 1.66 693.36 4.16 ;
      RECT  689.82 4.16 690.28 664.66 ;
      RECT  693.22 4.16 693.36 664.66 ;
      RECT  689.82 664.66 690.28 667.16 ;
      RECT  693.22 664.66 693.36 667.16 ;
   END
END    sky130_sram_4kbyte_1rw1r_32x1024_8
END    LIBRARY
