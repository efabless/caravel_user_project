magic
tech sky130A
magscale 1 2
timestamp 1617295513
<< obsli1 >>
rect 1104 833 118864 117521
<< obsm1 >>
rect 106 8 119862 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2318 119200 2374 120000
rect 3238 119200 3294 120000
rect 4158 119200 4214 120000
rect 5078 119200 5134 120000
rect 5998 119200 6054 120000
rect 6918 119200 6974 120000
rect 7838 119200 7894 120000
rect 8758 119200 8814 120000
rect 9770 119200 9826 120000
rect 10690 119200 10746 120000
rect 11610 119200 11666 120000
rect 12530 119200 12586 120000
rect 13450 119200 13506 120000
rect 14370 119200 14426 120000
rect 15290 119200 15346 120000
rect 16210 119200 16266 120000
rect 17130 119200 17186 120000
rect 18142 119200 18198 120000
rect 19062 119200 19118 120000
rect 19982 119200 20038 120000
rect 20902 119200 20958 120000
rect 21822 119200 21878 120000
rect 22742 119200 22798 120000
rect 23662 119200 23718 120000
rect 24582 119200 24638 120000
rect 25502 119200 25558 120000
rect 26514 119200 26570 120000
rect 27434 119200 27490 120000
rect 28354 119200 28410 120000
rect 29274 119200 29330 120000
rect 30194 119200 30250 120000
rect 31114 119200 31170 120000
rect 32034 119200 32090 120000
rect 32954 119200 33010 120000
rect 33874 119200 33930 120000
rect 34886 119200 34942 120000
rect 35806 119200 35862 120000
rect 36726 119200 36782 120000
rect 37646 119200 37702 120000
rect 38566 119200 38622 120000
rect 39486 119200 39542 120000
rect 40406 119200 40462 120000
rect 41326 119200 41382 120000
rect 42246 119200 42302 120000
rect 43166 119200 43222 120000
rect 44178 119200 44234 120000
rect 45098 119200 45154 120000
rect 46018 119200 46074 120000
rect 46938 119200 46994 120000
rect 47858 119200 47914 120000
rect 48778 119200 48834 120000
rect 49698 119200 49754 120000
rect 50618 119200 50674 120000
rect 51538 119200 51594 120000
rect 52550 119200 52606 120000
rect 53470 119200 53526 120000
rect 54390 119200 54446 120000
rect 55310 119200 55366 120000
rect 56230 119200 56286 120000
rect 57150 119200 57206 120000
rect 58070 119200 58126 120000
rect 58990 119200 59046 120000
rect 59910 119200 59966 120000
rect 60922 119200 60978 120000
rect 61842 119200 61898 120000
rect 62762 119200 62818 120000
rect 63682 119200 63738 120000
rect 64602 119200 64658 120000
rect 65522 119200 65578 120000
rect 66442 119200 66498 120000
rect 67362 119200 67418 120000
rect 68282 119200 68338 120000
rect 69294 119200 69350 120000
rect 70214 119200 70270 120000
rect 71134 119200 71190 120000
rect 72054 119200 72110 120000
rect 72974 119200 73030 120000
rect 73894 119200 73950 120000
rect 74814 119200 74870 120000
rect 75734 119200 75790 120000
rect 76654 119200 76710 120000
rect 77666 119200 77722 120000
rect 78586 119200 78642 120000
rect 79506 119200 79562 120000
rect 80426 119200 80482 120000
rect 81346 119200 81402 120000
rect 82266 119200 82322 120000
rect 83186 119200 83242 120000
rect 84106 119200 84162 120000
rect 85026 119200 85082 120000
rect 85946 119200 86002 120000
rect 86958 119200 87014 120000
rect 87878 119200 87934 120000
rect 88798 119200 88854 120000
rect 89718 119200 89774 120000
rect 90638 119200 90694 120000
rect 91558 119200 91614 120000
rect 92478 119200 92534 120000
rect 93398 119200 93454 120000
rect 94318 119200 94374 120000
rect 95330 119200 95386 120000
rect 96250 119200 96306 120000
rect 97170 119200 97226 120000
rect 98090 119200 98146 120000
rect 99010 119200 99066 120000
rect 99930 119200 99986 120000
rect 100850 119200 100906 120000
rect 101770 119200 101826 120000
rect 102690 119200 102746 120000
rect 103702 119200 103758 120000
rect 104622 119200 104678 120000
rect 105542 119200 105598 120000
rect 106462 119200 106518 120000
rect 107382 119200 107438 120000
rect 108302 119200 108358 120000
rect 109222 119200 109278 120000
rect 110142 119200 110198 120000
rect 111062 119200 111118 120000
rect 112074 119200 112130 120000
rect 112994 119200 113050 120000
rect 113914 119200 113970 120000
rect 114834 119200 114890 120000
rect 115754 119200 115810 120000
rect 116674 119200 116730 120000
rect 117594 119200 117650 120000
rect 118514 119200 118570 120000
rect 119434 119200 119490 120000
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1490 0 1546 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55402 0 55458 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62762 0 62818 800
rect 62946 0 63002 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69386 0 69442 800
rect 69570 0 69626 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70582 0 70638 800
rect 70858 0 70914 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72514 0 72570 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91834 0 91890 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 96986 0 97042 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98458 0 98514 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99194 0 99250 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101402 0 101458 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102138 0 102194 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106094 0 106150 800
rect 106278 0 106334 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109038 0 109094 800
rect 109222 0 109278 800
rect 109498 0 109554 800
rect 109774 0 109830 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110694 0 110750 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112166 0 112222 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113454 0 113510 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118054 0 118110 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119802 0 119858 800
<< obsm2 >>
rect 112 119144 422 119200
rect 590 119144 1342 119200
rect 1510 119144 2262 119200
rect 2430 119144 3182 119200
rect 3350 119144 4102 119200
rect 4270 119144 5022 119200
rect 5190 119144 5942 119200
rect 6110 119144 6862 119200
rect 7030 119144 7782 119200
rect 7950 119144 8702 119200
rect 8870 119144 9714 119200
rect 9882 119144 10634 119200
rect 10802 119144 11554 119200
rect 11722 119144 12474 119200
rect 12642 119144 13394 119200
rect 13562 119144 14314 119200
rect 14482 119144 15234 119200
rect 15402 119144 16154 119200
rect 16322 119144 17074 119200
rect 17242 119144 18086 119200
rect 18254 119144 19006 119200
rect 19174 119144 19926 119200
rect 20094 119144 20846 119200
rect 21014 119144 21766 119200
rect 21934 119144 22686 119200
rect 22854 119144 23606 119200
rect 23774 119144 24526 119200
rect 24694 119144 25446 119200
rect 25614 119144 26458 119200
rect 26626 119144 27378 119200
rect 27546 119144 28298 119200
rect 28466 119144 29218 119200
rect 29386 119144 30138 119200
rect 30306 119144 31058 119200
rect 31226 119144 31978 119200
rect 32146 119144 32898 119200
rect 33066 119144 33818 119200
rect 33986 119144 34830 119200
rect 34998 119144 35750 119200
rect 35918 119144 36670 119200
rect 36838 119144 37590 119200
rect 37758 119144 38510 119200
rect 38678 119144 39430 119200
rect 39598 119144 40350 119200
rect 40518 119144 41270 119200
rect 41438 119144 42190 119200
rect 42358 119144 43110 119200
rect 43278 119144 44122 119200
rect 44290 119144 45042 119200
rect 45210 119144 45962 119200
rect 46130 119144 46882 119200
rect 47050 119144 47802 119200
rect 47970 119144 48722 119200
rect 48890 119144 49642 119200
rect 49810 119144 50562 119200
rect 50730 119144 51482 119200
rect 51650 119144 52494 119200
rect 52662 119144 53414 119200
rect 53582 119144 54334 119200
rect 54502 119144 55254 119200
rect 55422 119144 56174 119200
rect 56342 119144 57094 119200
rect 57262 119144 58014 119200
rect 58182 119144 58934 119200
rect 59102 119144 59854 119200
rect 60022 119144 60866 119200
rect 61034 119144 61786 119200
rect 61954 119144 62706 119200
rect 62874 119144 63626 119200
rect 63794 119144 64546 119200
rect 64714 119144 65466 119200
rect 65634 119144 66386 119200
rect 66554 119144 67306 119200
rect 67474 119144 68226 119200
rect 68394 119144 69238 119200
rect 69406 119144 70158 119200
rect 70326 119144 71078 119200
rect 71246 119144 71998 119200
rect 72166 119144 72918 119200
rect 73086 119144 73838 119200
rect 74006 119144 74758 119200
rect 74926 119144 75678 119200
rect 75846 119144 76598 119200
rect 76766 119144 77610 119200
rect 77778 119144 78530 119200
rect 78698 119144 79450 119200
rect 79618 119144 80370 119200
rect 80538 119144 81290 119200
rect 81458 119144 82210 119200
rect 82378 119144 83130 119200
rect 83298 119144 84050 119200
rect 84218 119144 84970 119200
rect 85138 119144 85890 119200
rect 86058 119144 86902 119200
rect 87070 119144 87822 119200
rect 87990 119144 88742 119200
rect 88910 119144 89662 119200
rect 89830 119144 90582 119200
rect 90750 119144 91502 119200
rect 91670 119144 92422 119200
rect 92590 119144 93342 119200
rect 93510 119144 94262 119200
rect 94430 119144 95274 119200
rect 95442 119144 96194 119200
rect 96362 119144 97114 119200
rect 97282 119144 98034 119200
rect 98202 119144 98954 119200
rect 99122 119144 99874 119200
rect 100042 119144 100794 119200
rect 100962 119144 101714 119200
rect 101882 119144 102634 119200
rect 102802 119144 103646 119200
rect 103814 119144 104566 119200
rect 104734 119144 105486 119200
rect 105654 119144 106406 119200
rect 106574 119144 107326 119200
rect 107494 119144 108246 119200
rect 108414 119144 109166 119200
rect 109334 119144 110086 119200
rect 110254 119144 111006 119200
rect 111174 119144 112018 119200
rect 112186 119144 112938 119200
rect 113106 119144 113858 119200
rect 114026 119144 114778 119200
rect 114946 119144 115698 119200
rect 115866 119144 116618 119200
rect 116786 119144 117538 119200
rect 117706 119144 118458 119200
rect 118626 119144 119378 119200
rect 119546 119144 119856 119200
rect 112 856 119856 119144
rect 222 2 238 856
rect 406 2 514 856
rect 682 2 698 856
rect 866 2 974 856
rect 1142 2 1250 856
rect 1418 2 1434 856
rect 1602 2 1710 856
rect 1878 2 1986 856
rect 2154 2 2170 856
rect 2338 2 2446 856
rect 2614 2 2722 856
rect 2890 2 2906 856
rect 3074 2 3182 856
rect 3350 2 3458 856
rect 3626 2 3642 856
rect 3810 2 3918 856
rect 4086 2 4194 856
rect 4362 2 4378 856
rect 4546 2 4654 856
rect 4822 2 4930 856
rect 5098 2 5114 856
rect 5282 2 5390 856
rect 5558 2 5666 856
rect 5834 2 5850 856
rect 6018 2 6126 856
rect 6294 2 6402 856
rect 6570 2 6586 856
rect 6754 2 6862 856
rect 7030 2 7138 856
rect 7306 2 7322 856
rect 7490 2 7598 856
rect 7766 2 7874 856
rect 8042 2 8058 856
rect 8226 2 8334 856
rect 8502 2 8610 856
rect 8778 2 8794 856
rect 8962 2 9070 856
rect 9238 2 9346 856
rect 9514 2 9530 856
rect 9698 2 9806 856
rect 9974 2 10082 856
rect 10250 2 10266 856
rect 10434 2 10542 856
rect 10710 2 10818 856
rect 10986 2 11002 856
rect 11170 2 11278 856
rect 11446 2 11554 856
rect 11722 2 11738 856
rect 11906 2 12014 856
rect 12182 2 12290 856
rect 12458 2 12474 856
rect 12642 2 12750 856
rect 12918 2 13026 856
rect 13194 2 13210 856
rect 13378 2 13486 856
rect 13654 2 13762 856
rect 13930 2 13946 856
rect 14114 2 14222 856
rect 14390 2 14498 856
rect 14666 2 14682 856
rect 14850 2 14958 856
rect 15126 2 15142 856
rect 15310 2 15418 856
rect 15586 2 15694 856
rect 15862 2 15878 856
rect 16046 2 16154 856
rect 16322 2 16430 856
rect 16598 2 16614 856
rect 16782 2 16890 856
rect 17058 2 17166 856
rect 17334 2 17350 856
rect 17518 2 17626 856
rect 17794 2 17902 856
rect 18070 2 18086 856
rect 18254 2 18362 856
rect 18530 2 18638 856
rect 18806 2 18822 856
rect 18990 2 19098 856
rect 19266 2 19374 856
rect 19542 2 19558 856
rect 19726 2 19834 856
rect 20002 2 20110 856
rect 20278 2 20294 856
rect 20462 2 20570 856
rect 20738 2 20846 856
rect 21014 2 21030 856
rect 21198 2 21306 856
rect 21474 2 21582 856
rect 21750 2 21766 856
rect 21934 2 22042 856
rect 22210 2 22318 856
rect 22486 2 22502 856
rect 22670 2 22778 856
rect 22946 2 23054 856
rect 23222 2 23238 856
rect 23406 2 23514 856
rect 23682 2 23790 856
rect 23958 2 23974 856
rect 24142 2 24250 856
rect 24418 2 24526 856
rect 24694 2 24710 856
rect 24878 2 24986 856
rect 25154 2 25262 856
rect 25430 2 25446 856
rect 25614 2 25722 856
rect 25890 2 25998 856
rect 26166 2 26182 856
rect 26350 2 26458 856
rect 26626 2 26734 856
rect 26902 2 26918 856
rect 27086 2 27194 856
rect 27362 2 27470 856
rect 27638 2 27654 856
rect 27822 2 27930 856
rect 28098 2 28206 856
rect 28374 2 28390 856
rect 28558 2 28666 856
rect 28834 2 28942 856
rect 29110 2 29126 856
rect 29294 2 29402 856
rect 29570 2 29678 856
rect 29846 2 29862 856
rect 30030 2 30138 856
rect 30306 2 30322 856
rect 30490 2 30598 856
rect 30766 2 30874 856
rect 31042 2 31058 856
rect 31226 2 31334 856
rect 31502 2 31610 856
rect 31778 2 31794 856
rect 31962 2 32070 856
rect 32238 2 32346 856
rect 32514 2 32530 856
rect 32698 2 32806 856
rect 32974 2 33082 856
rect 33250 2 33266 856
rect 33434 2 33542 856
rect 33710 2 33818 856
rect 33986 2 34002 856
rect 34170 2 34278 856
rect 34446 2 34554 856
rect 34722 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35290 856
rect 35458 2 35474 856
rect 35642 2 35750 856
rect 35918 2 36026 856
rect 36194 2 36210 856
rect 36378 2 36486 856
rect 36654 2 36762 856
rect 36930 2 36946 856
rect 37114 2 37222 856
rect 37390 2 37498 856
rect 37666 2 37682 856
rect 37850 2 37958 856
rect 38126 2 38234 856
rect 38402 2 38418 856
rect 38586 2 38694 856
rect 38862 2 38970 856
rect 39138 2 39154 856
rect 39322 2 39430 856
rect 39598 2 39706 856
rect 39874 2 39890 856
rect 40058 2 40166 856
rect 40334 2 40442 856
rect 40610 2 40626 856
rect 40794 2 40902 856
rect 41070 2 41178 856
rect 41346 2 41362 856
rect 41530 2 41638 856
rect 41806 2 41914 856
rect 42082 2 42098 856
rect 42266 2 42374 856
rect 42542 2 42650 856
rect 42818 2 42834 856
rect 43002 2 43110 856
rect 43278 2 43386 856
rect 43554 2 43570 856
rect 43738 2 43846 856
rect 44014 2 44122 856
rect 44290 2 44306 856
rect 44474 2 44582 856
rect 44750 2 44858 856
rect 45026 2 45042 856
rect 45210 2 45318 856
rect 45486 2 45502 856
rect 45670 2 45778 856
rect 45946 2 46054 856
rect 46222 2 46238 856
rect 46406 2 46514 856
rect 46682 2 46790 856
rect 46958 2 46974 856
rect 47142 2 47250 856
rect 47418 2 47526 856
rect 47694 2 47710 856
rect 47878 2 47986 856
rect 48154 2 48262 856
rect 48430 2 48446 856
rect 48614 2 48722 856
rect 48890 2 48998 856
rect 49166 2 49182 856
rect 49350 2 49458 856
rect 49626 2 49734 856
rect 49902 2 49918 856
rect 50086 2 50194 856
rect 50362 2 50470 856
rect 50638 2 50654 856
rect 50822 2 50930 856
rect 51098 2 51206 856
rect 51374 2 51390 856
rect 51558 2 51666 856
rect 51834 2 51942 856
rect 52110 2 52126 856
rect 52294 2 52402 856
rect 52570 2 52678 856
rect 52846 2 52862 856
rect 53030 2 53138 856
rect 53306 2 53414 856
rect 53582 2 53598 856
rect 53766 2 53874 856
rect 54042 2 54150 856
rect 54318 2 54334 856
rect 54502 2 54610 856
rect 54778 2 54886 856
rect 55054 2 55070 856
rect 55238 2 55346 856
rect 55514 2 55622 856
rect 55790 2 55806 856
rect 55974 2 56082 856
rect 56250 2 56358 856
rect 56526 2 56542 856
rect 56710 2 56818 856
rect 56986 2 57094 856
rect 57262 2 57278 856
rect 57446 2 57554 856
rect 57722 2 57830 856
rect 57998 2 58014 856
rect 58182 2 58290 856
rect 58458 2 58566 856
rect 58734 2 58750 856
rect 58918 2 59026 856
rect 59194 2 59302 856
rect 59470 2 59486 856
rect 59654 2 59762 856
rect 59930 2 60038 856
rect 60206 2 60222 856
rect 60390 2 60498 856
rect 60666 2 60682 856
rect 60850 2 60958 856
rect 61126 2 61234 856
rect 61402 2 61418 856
rect 61586 2 61694 856
rect 61862 2 61970 856
rect 62138 2 62154 856
rect 62322 2 62430 856
rect 62598 2 62706 856
rect 62874 2 62890 856
rect 63058 2 63166 856
rect 63334 2 63442 856
rect 63610 2 63626 856
rect 63794 2 63902 856
rect 64070 2 64178 856
rect 64346 2 64362 856
rect 64530 2 64638 856
rect 64806 2 64914 856
rect 65082 2 65098 856
rect 65266 2 65374 856
rect 65542 2 65650 856
rect 65818 2 65834 856
rect 66002 2 66110 856
rect 66278 2 66386 856
rect 66554 2 66570 856
rect 66738 2 66846 856
rect 67014 2 67122 856
rect 67290 2 67306 856
rect 67474 2 67582 856
rect 67750 2 67858 856
rect 68026 2 68042 856
rect 68210 2 68318 856
rect 68486 2 68594 856
rect 68762 2 68778 856
rect 68946 2 69054 856
rect 69222 2 69330 856
rect 69498 2 69514 856
rect 69682 2 69790 856
rect 69958 2 70066 856
rect 70234 2 70250 856
rect 70418 2 70526 856
rect 70694 2 70802 856
rect 70970 2 70986 856
rect 71154 2 71262 856
rect 71430 2 71538 856
rect 71706 2 71722 856
rect 71890 2 71998 856
rect 72166 2 72274 856
rect 72442 2 72458 856
rect 72626 2 72734 856
rect 72902 2 73010 856
rect 73178 2 73194 856
rect 73362 2 73470 856
rect 73638 2 73746 856
rect 73914 2 73930 856
rect 74098 2 74206 856
rect 74374 2 74482 856
rect 74650 2 74666 856
rect 74834 2 74942 856
rect 75110 2 75126 856
rect 75294 2 75402 856
rect 75570 2 75678 856
rect 75846 2 75862 856
rect 76030 2 76138 856
rect 76306 2 76414 856
rect 76582 2 76598 856
rect 76766 2 76874 856
rect 77042 2 77150 856
rect 77318 2 77334 856
rect 77502 2 77610 856
rect 77778 2 77886 856
rect 78054 2 78070 856
rect 78238 2 78346 856
rect 78514 2 78622 856
rect 78790 2 78806 856
rect 78974 2 79082 856
rect 79250 2 79358 856
rect 79526 2 79542 856
rect 79710 2 79818 856
rect 79986 2 80094 856
rect 80262 2 80278 856
rect 80446 2 80554 856
rect 80722 2 80830 856
rect 80998 2 81014 856
rect 81182 2 81290 856
rect 81458 2 81566 856
rect 81734 2 81750 856
rect 81918 2 82026 856
rect 82194 2 82302 856
rect 82470 2 82486 856
rect 82654 2 82762 856
rect 82930 2 83038 856
rect 83206 2 83222 856
rect 83390 2 83498 856
rect 83666 2 83774 856
rect 83942 2 83958 856
rect 84126 2 84234 856
rect 84402 2 84510 856
rect 84678 2 84694 856
rect 84862 2 84970 856
rect 85138 2 85246 856
rect 85414 2 85430 856
rect 85598 2 85706 856
rect 85874 2 85982 856
rect 86150 2 86166 856
rect 86334 2 86442 856
rect 86610 2 86718 856
rect 86886 2 86902 856
rect 87070 2 87178 856
rect 87346 2 87454 856
rect 87622 2 87638 856
rect 87806 2 87914 856
rect 88082 2 88190 856
rect 88358 2 88374 856
rect 88542 2 88650 856
rect 88818 2 88926 856
rect 89094 2 89110 856
rect 89278 2 89386 856
rect 89554 2 89662 856
rect 89830 2 89846 856
rect 90014 2 90122 856
rect 90290 2 90306 856
rect 90474 2 90582 856
rect 90750 2 90858 856
rect 91026 2 91042 856
rect 91210 2 91318 856
rect 91486 2 91594 856
rect 91762 2 91778 856
rect 91946 2 92054 856
rect 92222 2 92330 856
rect 92498 2 92514 856
rect 92682 2 92790 856
rect 92958 2 93066 856
rect 93234 2 93250 856
rect 93418 2 93526 856
rect 93694 2 93802 856
rect 93970 2 93986 856
rect 94154 2 94262 856
rect 94430 2 94538 856
rect 94706 2 94722 856
rect 94890 2 94998 856
rect 95166 2 95274 856
rect 95442 2 95458 856
rect 95626 2 95734 856
rect 95902 2 96010 856
rect 96178 2 96194 856
rect 96362 2 96470 856
rect 96638 2 96746 856
rect 96914 2 96930 856
rect 97098 2 97206 856
rect 97374 2 97482 856
rect 97650 2 97666 856
rect 97834 2 97942 856
rect 98110 2 98218 856
rect 98386 2 98402 856
rect 98570 2 98678 856
rect 98846 2 98954 856
rect 99122 2 99138 856
rect 99306 2 99414 856
rect 99582 2 99690 856
rect 99858 2 99874 856
rect 100042 2 100150 856
rect 100318 2 100426 856
rect 100594 2 100610 856
rect 100778 2 100886 856
rect 101054 2 101162 856
rect 101330 2 101346 856
rect 101514 2 101622 856
rect 101790 2 101898 856
rect 102066 2 102082 856
rect 102250 2 102358 856
rect 102526 2 102634 856
rect 102802 2 102818 856
rect 102986 2 103094 856
rect 103262 2 103370 856
rect 103538 2 103554 856
rect 103722 2 103830 856
rect 103998 2 104106 856
rect 104274 2 104290 856
rect 104458 2 104566 856
rect 104734 2 104842 856
rect 105010 2 105026 856
rect 105194 2 105302 856
rect 105470 2 105486 856
rect 105654 2 105762 856
rect 105930 2 106038 856
rect 106206 2 106222 856
rect 106390 2 106498 856
rect 106666 2 106774 856
rect 106942 2 106958 856
rect 107126 2 107234 856
rect 107402 2 107510 856
rect 107678 2 107694 856
rect 107862 2 107970 856
rect 108138 2 108246 856
rect 108414 2 108430 856
rect 108598 2 108706 856
rect 108874 2 108982 856
rect 109150 2 109166 856
rect 109334 2 109442 856
rect 109610 2 109718 856
rect 109886 2 109902 856
rect 110070 2 110178 856
rect 110346 2 110454 856
rect 110622 2 110638 856
rect 110806 2 110914 856
rect 111082 2 111190 856
rect 111358 2 111374 856
rect 111542 2 111650 856
rect 111818 2 111926 856
rect 112094 2 112110 856
rect 112278 2 112386 856
rect 112554 2 112662 856
rect 112830 2 112846 856
rect 113014 2 113122 856
rect 113290 2 113398 856
rect 113566 2 113582 856
rect 113750 2 113858 856
rect 114026 2 114134 856
rect 114302 2 114318 856
rect 114486 2 114594 856
rect 114762 2 114870 856
rect 115038 2 115054 856
rect 115222 2 115330 856
rect 115498 2 115606 856
rect 115774 2 115790 856
rect 115958 2 116066 856
rect 116234 2 116342 856
rect 116510 2 116526 856
rect 116694 2 116802 856
rect 116970 2 117078 856
rect 117246 2 117262 856
rect 117430 2 117538 856
rect 117706 2 117814 856
rect 117982 2 117998 856
rect 118166 2 118274 856
rect 118442 2 118550 856
rect 118718 2 118734 856
rect 118902 2 119010 856
rect 119178 2 119286 856
rect 119454 2 119470 856
rect 119638 2 119746 856
<< obsm3 >>
rect 2681 716 112048 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
<< obsm4 >>
rect 7971 2048 19488 13837
rect 19968 2096 20148 13837
rect 20628 2096 20808 13837
rect 21288 2096 21468 13837
rect 21948 2096 34848 13837
rect 19968 2048 34848 2096
rect 35328 2096 35508 13837
rect 35988 2096 36168 13837
rect 36648 2096 36828 13837
rect 37308 2096 50208 13837
rect 35328 2048 50208 2096
rect 50688 2096 50868 13837
rect 51348 2096 51528 13837
rect 52008 2096 52188 13837
rect 52668 2096 65445 13837
rect 50688 2048 65445 2096
rect 7971 715 65445 2048
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 28354 119200 28410 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 31114 119200 31170 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 33874 119200 33930 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 36726 119200 36782 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 39486 119200 39542 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 42246 119200 42302 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 45098 119200 45154 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 47858 119200 47914 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 50618 119200 50674 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 53470 119200 53526 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3238 119200 3294 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 56230 119200 56286 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 58990 119200 59046 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 61842 119200 61898 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 64602 119200 64658 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 67362 119200 67418 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 70214 119200 70270 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 72974 119200 73030 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 75734 119200 75790 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 78586 119200 78642 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 81346 119200 81402 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5998 119200 6054 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 84106 119200 84162 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 86958 119200 87014 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 89718 119200 89774 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 92478 119200 92534 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 95330 119200 95386 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 98090 119200 98146 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 100850 119200 100906 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 103702 119200 103758 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 106462 119200 106518 120000 6 io_in[38]
port 32 nsew signal input
rlabel metal2 s 109222 119200 109278 120000 6 io_in[39]
port 33 nsew signal input
rlabel metal2 s 8758 119200 8814 120000 6 io_in[3]
port 34 nsew signal input
rlabel metal2 s 112074 119200 112130 120000 6 io_in[40]
port 35 nsew signal input
rlabel metal2 s 114834 119200 114890 120000 6 io_in[41]
port 36 nsew signal input
rlabel metal2 s 117594 119200 117650 120000 6 io_in[42]
port 37 nsew signal input
rlabel metal2 s 11610 119200 11666 120000 6 io_in[4]
port 38 nsew signal input
rlabel metal2 s 14370 119200 14426 120000 6 io_in[5]
port 39 nsew signal input
rlabel metal2 s 17130 119200 17186 120000 6 io_in[6]
port 40 nsew signal input
rlabel metal2 s 19982 119200 20038 120000 6 io_in[7]
port 41 nsew signal input
rlabel metal2 s 22742 119200 22798 120000 6 io_in[8]
port 42 nsew signal input
rlabel metal2 s 25502 119200 25558 120000 6 io_in[9]
port 43 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 io_oeb[0]
port 44 nsew signal output
rlabel metal2 s 29274 119200 29330 120000 6 io_oeb[10]
port 45 nsew signal output
rlabel metal2 s 32034 119200 32090 120000 6 io_oeb[11]
port 46 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_oeb[12]
port 47 nsew signal output
rlabel metal2 s 37646 119200 37702 120000 6 io_oeb[13]
port 48 nsew signal output
rlabel metal2 s 40406 119200 40462 120000 6 io_oeb[14]
port 49 nsew signal output
rlabel metal2 s 43166 119200 43222 120000 6 io_oeb[15]
port 50 nsew signal output
rlabel metal2 s 46018 119200 46074 120000 6 io_oeb[16]
port 51 nsew signal output
rlabel metal2 s 48778 119200 48834 120000 6 io_oeb[17]
port 52 nsew signal output
rlabel metal2 s 51538 119200 51594 120000 6 io_oeb[18]
port 53 nsew signal output
rlabel metal2 s 54390 119200 54446 120000 6 io_oeb[19]
port 54 nsew signal output
rlabel metal2 s 4158 119200 4214 120000 6 io_oeb[1]
port 55 nsew signal output
rlabel metal2 s 57150 119200 57206 120000 6 io_oeb[20]
port 56 nsew signal output
rlabel metal2 s 59910 119200 59966 120000 6 io_oeb[21]
port 57 nsew signal output
rlabel metal2 s 62762 119200 62818 120000 6 io_oeb[22]
port 58 nsew signal output
rlabel metal2 s 65522 119200 65578 120000 6 io_oeb[23]
port 59 nsew signal output
rlabel metal2 s 68282 119200 68338 120000 6 io_oeb[24]
port 60 nsew signal output
rlabel metal2 s 71134 119200 71190 120000 6 io_oeb[25]
port 61 nsew signal output
rlabel metal2 s 73894 119200 73950 120000 6 io_oeb[26]
port 62 nsew signal output
rlabel metal2 s 76654 119200 76710 120000 6 io_oeb[27]
port 63 nsew signal output
rlabel metal2 s 79506 119200 79562 120000 6 io_oeb[28]
port 64 nsew signal output
rlabel metal2 s 82266 119200 82322 120000 6 io_oeb[29]
port 65 nsew signal output
rlabel metal2 s 6918 119200 6974 120000 6 io_oeb[2]
port 66 nsew signal output
rlabel metal2 s 85026 119200 85082 120000 6 io_oeb[30]
port 67 nsew signal output
rlabel metal2 s 87878 119200 87934 120000 6 io_oeb[31]
port 68 nsew signal output
rlabel metal2 s 90638 119200 90694 120000 6 io_oeb[32]
port 69 nsew signal output
rlabel metal2 s 93398 119200 93454 120000 6 io_oeb[33]
port 70 nsew signal output
rlabel metal2 s 96250 119200 96306 120000 6 io_oeb[34]
port 71 nsew signal output
rlabel metal2 s 99010 119200 99066 120000 6 io_oeb[35]
port 72 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 io_oeb[36]
port 73 nsew signal output
rlabel metal2 s 104622 119200 104678 120000 6 io_oeb[37]
port 74 nsew signal output
rlabel metal2 s 107382 119200 107438 120000 6 io_oeb[38]
port 75 nsew signal output
rlabel metal2 s 110142 119200 110198 120000 6 io_oeb[39]
port 76 nsew signal output
rlabel metal2 s 9770 119200 9826 120000 6 io_oeb[3]
port 77 nsew signal output
rlabel metal2 s 112994 119200 113050 120000 6 io_oeb[40]
port 78 nsew signal output
rlabel metal2 s 115754 119200 115810 120000 6 io_oeb[41]
port 79 nsew signal output
rlabel metal2 s 118514 119200 118570 120000 6 io_oeb[42]
port 80 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 15290 119200 15346 120000 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 18142 119200 18198 120000 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 20902 119200 20958 120000 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 23662 119200 23718 120000 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 26514 119200 26570 120000 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 2318 119200 2374 120000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 30194 119200 30250 120000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 32954 119200 33010 120000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 35806 119200 35862 120000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 38566 119200 38622 120000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 41326 119200 41382 120000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 44178 119200 44234 120000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 49698 119200 49754 120000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 52550 119200 52606 120000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 55310 119200 55366 120000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 5078 119200 5134 120000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 58070 119200 58126 120000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 60922 119200 60978 120000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 63682 119200 63738 120000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 66442 119200 66498 120000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 69294 119200 69350 120000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 72054 119200 72110 120000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 74814 119200 74870 120000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 77666 119200 77722 120000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 80426 119200 80482 120000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 83186 119200 83242 120000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 85946 119200 86002 120000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 88798 119200 88854 120000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 91558 119200 91614 120000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 94318 119200 94374 120000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 97170 119200 97226 120000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 99930 119200 99986 120000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 102690 119200 102746 120000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 105542 119200 105598 120000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 108302 119200 108358 120000 6 io_out[38]
port 118 nsew signal output
rlabel metal2 s 111062 119200 111118 120000 6 io_out[39]
port 119 nsew signal output
rlabel metal2 s 10690 119200 10746 120000 6 io_out[3]
port 120 nsew signal output
rlabel metal2 s 113914 119200 113970 120000 6 io_out[40]
port 121 nsew signal output
rlabel metal2 s 116674 119200 116730 120000 6 io_out[41]
port 122 nsew signal output
rlabel metal2 s 119434 119200 119490 120000 6 io_out[42]
port 123 nsew signal output
rlabel metal2 s 13450 119200 13506 120000 6 io_out[4]
port 124 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 io_out[5]
port 125 nsew signal output
rlabel metal2 s 19062 119200 19118 120000 6 io_out[6]
port 126 nsew signal output
rlabel metal2 s 21822 119200 21878 120000 6 io_out[7]
port 127 nsew signal output
rlabel metal2 s 24582 119200 24638 120000 6 io_out[8]
port 128 nsew signal output
rlabel metal2 s 27434 119200 27490 120000 6 io_out[9]
port 129 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 la_data_in[0]
port 130 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[100]
port 131 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[101]
port 132 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[102]
port 133 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[103]
port 134 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[104]
port 135 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[105]
port 136 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[106]
port 137 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[107]
port 138 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[108]
port 139 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[109]
port 140 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[10]
port 141 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[110]
port 142 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[111]
port 143 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[112]
port 144 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[113]
port 145 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[114]
port 146 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[115]
port 147 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[116]
port 148 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[117]
port 149 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[118]
port 150 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[119]
port 151 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_data_in[11]
port 152 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[120]
port 153 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[121]
port 154 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[122]
port 155 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[123]
port 156 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[124]
port 157 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[125]
port 158 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[126]
port 159 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[127]
port 160 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[12]
port 161 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_data_in[13]
port 162 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[14]
port 163 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[15]
port 164 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_in[16]
port 165 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_in[17]
port 166 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[18]
port 167 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[19]
port 168 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[1]
port 169 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[20]
port 170 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[21]
port 171 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[22]
port 172 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[23]
port 173 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[24]
port 174 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[25]
port 175 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[26]
port 176 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[27]
port 177 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[28]
port 178 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[29]
port 179 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_data_in[2]
port 180 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[30]
port 181 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[31]
port 182 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[32]
port 183 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[33]
port 184 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[34]
port 185 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[35]
port 186 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[36]
port 187 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[37]
port 188 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[38]
port 189 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[39]
port 190 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[3]
port 191 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[40]
port 192 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[41]
port 193 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[42]
port 194 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[43]
port 195 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[44]
port 196 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[45]
port 197 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[46]
port 198 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[47]
port 199 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[48]
port 200 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[49]
port 201 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[4]
port 202 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[50]
port 203 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[51]
port 204 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[52]
port 205 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[53]
port 206 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[54]
port 207 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[55]
port 208 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_data_in[56]
port 209 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[57]
port 210 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[58]
port 211 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[59]
port 212 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[5]
port 213 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[60]
port 214 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[61]
port 215 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[62]
port 216 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[63]
port 217 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[64]
port 218 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[65]
port 219 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[66]
port 220 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[67]
port 221 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[68]
port 222 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[69]
port 223 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[6]
port 224 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[70]
port 225 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[71]
port 226 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[72]
port 227 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[73]
port 228 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[74]
port 229 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[75]
port 230 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[76]
port 231 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[77]
port 232 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[78]
port 233 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[79]
port 234 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_data_in[7]
port 235 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[80]
port 236 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[81]
port 237 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[82]
port 238 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[83]
port 239 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[84]
port 240 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[85]
port 241 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[86]
port 242 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[87]
port 243 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[88]
port 244 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[89]
port 245 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[8]
port 246 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[90]
port 247 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[91]
port 248 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[92]
port 249 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[93]
port 250 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_data_in[94]
port 251 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[95]
port 252 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[96]
port 253 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[97]
port 254 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[98]
port 255 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[99]
port 256 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[9]
port 257 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_out[0]
port 258 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[100]
port 259 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[101]
port 260 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[102]
port 261 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[103]
port 262 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 la_data_out[104]
port 263 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[105]
port 264 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[106]
port 265 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[107]
port 266 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[108]
port 267 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 la_data_out[109]
port 268 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 la_data_out[10]
port 269 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[110]
port 270 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[111]
port 271 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[112]
port 272 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[113]
port 273 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_data_out[114]
port 274 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[115]
port 275 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[116]
port 276 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[117]
port 277 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[118]
port 278 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[119]
port 279 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 la_data_out[11]
port 280 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[120]
port 281 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[121]
port 282 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[122]
port 283 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[123]
port 284 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[124]
port 285 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[125]
port 286 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[126]
port 287 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[127]
port 288 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[12]
port 289 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[13]
port 290 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[14]
port 291 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[15]
port 292 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[16]
port 293 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[17]
port 294 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[18]
port 295 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[19]
port 296 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 la_data_out[1]
port 297 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[20]
port 298 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[21]
port 299 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[22]
port 300 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[23]
port 301 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[24]
port 302 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[25]
port 303 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[26]
port 304 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[27]
port 305 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[28]
port 306 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[29]
port 307 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[2]
port 308 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[30]
port 309 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[31]
port 310 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[32]
port 311 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[33]
port 312 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[34]
port 313 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[35]
port 314 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[36]
port 315 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[37]
port 316 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[38]
port 317 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[39]
port 318 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 la_data_out[3]
port 319 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[40]
port 320 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[41]
port 321 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[42]
port 322 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[43]
port 323 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[44]
port 324 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[45]
port 325 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[46]
port 326 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[47]
port 327 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[48]
port 328 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[49]
port 329 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[4]
port 330 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[50]
port 331 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[51]
port 332 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[52]
port 333 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[53]
port 334 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[54]
port 335 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[55]
port 336 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 la_data_out[56]
port 337 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[57]
port 338 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[58]
port 339 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[59]
port 340 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 la_data_out[5]
port 341 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[60]
port 342 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[61]
port 343 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[62]
port 344 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[63]
port 345 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[64]
port 346 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[65]
port 347 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[66]
port 348 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[67]
port 349 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[68]
port 350 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[69]
port 351 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_data_out[6]
port 352 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[70]
port 353 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[71]
port 354 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[72]
port 355 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[73]
port 356 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[74]
port 357 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[75]
port 358 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[76]
port 359 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[77]
port 360 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[78]
port 361 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[79]
port 362 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[7]
port 363 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[80]
port 364 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[81]
port 365 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[82]
port 366 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[83]
port 367 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[84]
port 368 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 la_data_out[85]
port 369 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[86]
port 370 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[87]
port 371 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[88]
port 372 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[89]
port 373 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[8]
port 374 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[90]
port 375 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[91]
port 376 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[92]
port 377 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[93]
port 378 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[94]
port 379 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[95]
port 380 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[96]
port 381 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[97]
port 382 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[98]
port 383 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[99]
port 384 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[9]
port 385 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_oen[0]
port 386 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oen[100]
port 387 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oen[101]
port 388 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oen[102]
port 389 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_oen[103]
port 390 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oen[104]
port 391 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_oen[105]
port 392 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oen[106]
port 393 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oen[107]
port 394 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oen[108]
port 395 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oen[109]
port 396 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oen[10]
port 397 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oen[110]
port 398 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_oen[111]
port 399 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oen[112]
port 400 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_oen[113]
port 401 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oen[114]
port 402 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_oen[115]
port 403 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_oen[116]
port 404 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oen[117]
port 405 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oen[118]
port 406 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oen[119]
port 407 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 la_oen[11]
port 408 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oen[120]
port 409 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oen[121]
port 410 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_oen[122]
port 411 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oen[123]
port 412 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oen[124]
port 413 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_oen[125]
port 414 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oen[126]
port 415 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oen[127]
port 416 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_oen[12]
port 417 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oen[13]
port 418 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oen[14]
port 419 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oen[15]
port 420 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oen[16]
port 421 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oen[17]
port 422 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oen[18]
port 423 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oen[19]
port 424 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oen[1]
port 425 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oen[20]
port 426 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oen[21]
port 427 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oen[22]
port 428 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oen[23]
port 429 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oen[24]
port 430 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oen[25]
port 431 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oen[26]
port 432 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oen[27]
port 433 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oen[28]
port 434 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oen[29]
port 435 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_oen[2]
port 436 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oen[30]
port 437 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oen[31]
port 438 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oen[32]
port 439 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oen[33]
port 440 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oen[34]
port 441 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oen[35]
port 442 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oen[36]
port 443 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oen[37]
port 444 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oen[38]
port 445 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oen[39]
port 446 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oen[3]
port 447 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oen[40]
port 448 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oen[41]
port 449 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oen[42]
port 450 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oen[43]
port 451 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oen[44]
port 452 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oen[45]
port 453 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oen[46]
port 454 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oen[47]
port 455 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oen[48]
port 456 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oen[49]
port 457 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_oen[4]
port 458 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oen[50]
port 459 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oen[51]
port 460 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oen[52]
port 461 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oen[53]
port 462 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oen[54]
port 463 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oen[55]
port 464 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oen[56]
port 465 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oen[57]
port 466 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oen[58]
port 467 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oen[59]
port 468 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_oen[5]
port 469 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oen[60]
port 470 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oen[61]
port 471 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oen[62]
port 472 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oen[63]
port 473 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oen[64]
port 474 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oen[65]
port 475 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oen[66]
port 476 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oen[67]
port 477 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oen[68]
port 478 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oen[69]
port 479 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_oen[6]
port 480 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oen[70]
port 481 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oen[71]
port 482 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oen[72]
port 483 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oen[73]
port 484 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oen[74]
port 485 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oen[75]
port 486 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oen[76]
port 487 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oen[77]
port 488 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oen[78]
port 489 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oen[79]
port 490 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oen[7]
port 491 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oen[80]
port 492 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oen[81]
port 493 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oen[82]
port 494 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oen[83]
port 495 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oen[84]
port 496 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oen[85]
port 497 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oen[86]
port 498 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oen[87]
port 499 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oen[88]
port 500 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oen[89]
port 501 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oen[8]
port 502 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oen[90]
port 503 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oen[91]
port 504 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oen[92]
port 505 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oen[93]
port 506 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oen[94]
port 507 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oen[95]
port 508 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oen[96]
port 509 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oen[97]
port 510 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oen[98]
port 511 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oen[99]
port 512 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oen[9]
port 513 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 514 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 515 nsew signal input
rlabel metal2 s 570 0 626 800 6 wbs_ack_o
port 516 nsew signal output
rlabel metal2 s 1490 0 1546 800 6 wbs_adr_i[0]
port 517 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[10]
port 518 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[11]
port 519 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[12]
port 520 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[13]
port 521 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[14]
port 522 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[15]
port 523 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[16]
port 524 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[17]
port 525 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[18]
port 526 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[19]
port 527 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[1]
port 528 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[20]
port 529 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[21]
port 530 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[22]
port 531 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_adr_i[23]
port 532 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[24]
port 533 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[25]
port 534 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[26]
port 535 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[27]
port 536 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[28]
port 537 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[29]
port 538 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_adr_i[2]
port 539 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[30]
port 540 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[31]
port 541 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[3]
port 542 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[4]
port 543 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[5]
port 544 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[6]
port 545 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_adr_i[7]
port 546 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[8]
port 547 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[9]
port 548 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 549 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_i[0]
port 550 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[10]
port 551 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[11]
port 552 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[12]
port 553 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[13]
port 554 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[14]
port 555 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[15]
port 556 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[16]
port 557 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_i[17]
port 558 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[18]
port 559 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[19]
port 560 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_i[1]
port 561 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_i[20]
port 562 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[21]
port 563 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[22]
port 564 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[23]
port 565 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[24]
port 566 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[25]
port 567 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[26]
port 568 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[27]
port 569 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[28]
port 570 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[29]
port 571 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[2]
port 572 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[30]
port 573 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[31]
port 574 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_i[3]
port 575 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[4]
port 576 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[5]
port 577 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[6]
port 578 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[7]
port 579 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[8]
port 580 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[9]
port 581 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_o[0]
port 582 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[10]
port 583 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[11]
port 584 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[12]
port 585 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[13]
port 586 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_o[14]
port 587 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[15]
port 588 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[16]
port 589 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[17]
port 590 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[18]
port 591 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[19]
port 592 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[1]
port 593 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_o[20]
port 594 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[21]
port 595 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[22]
port 596 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[23]
port 597 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[24]
port 598 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[25]
port 599 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[26]
port 600 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[27]
port 601 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_o[28]
port 602 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[29]
port 603 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[2]
port 604 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[30]
port 605 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[31]
port 606 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_o[3]
port 607 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[4]
port 608 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[5]
port 609 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[6]
port 610 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[7]
port 611 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[8]
port 612 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[9]
port 613 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[0]
port 614 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[1]
port 615 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[2]
port 616 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[3]
port 617 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_stb_i
port 618 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_we_i
port 619 nsew signal input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 620 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 621 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 622 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 633 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 638 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 639 nsew power bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 640 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 644 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 645 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 646 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 648 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 649 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 650 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 651 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 120000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 6085594
string GDS_START 267896
<< end >>

